// This is the unpowered netlist.
module tiny_user_project (io_in,
    io_oeb,
    io_out);
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire net53;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net54;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net55;
 wire net83;
 wire net84;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net22;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net23;
 wire net42;
 wire net43;
 wire net44;
 wire net24;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire \mod.flipflop1.d ;
 wire \mod.flipflop1.q ;
 wire \mod.flipflop10.d ;
 wire \mod.flipflop11.d ;
 wire \mod.flipflop11.q ;
 wire \mod.flipflop12.d ;
 wire \mod.flipflop12.q ;
 wire \mod.flipflop13.q ;
 wire \mod.flipflop14.q ;
 wire \mod.flipflop15.d ;
 wire \mod.flipflop16.d ;
 wire \mod.flipflop17.d ;
 wire \mod.flipflop18.d ;
 wire \mod.flipflop18.q ;
 wire \mod.flipflop19.q ;
 wire \mod.flipflop2.d ;
 wire \mod.flipflop2.q ;
 wire \mod.flipflop20.q ;
 wire \mod.flipflop21.d ;
 wire \mod.flipflop21.q ;
 wire \mod.flipflop22.q ;
 wire \mod.flipflop23.q ;
 wire \mod.flipflop24.q ;
 wire \mod.flipflop25.q ;
 wire \mod.flipflop26.q ;
 wire \mod.flipflop27.d ;
 wire \mod.flipflop27.q ;
 wire \mod.flipflop28.q ;
 wire \mod.flipflop29.d ;
 wire \mod.flipflop29.q ;
 wire \mod.flipflop3.q ;
 wire \mod.flipflop30.q ;
 wire \mod.flipflop31.q ;
 wire \mod.flipflop32.d ;
 wire \mod.flipflop32.q ;
 wire \mod.flipflop33.d ;
 wire \mod.flipflop33.q ;
 wire \mod.flipflop34.d ;
 wire \mod.flipflop34.q ;
 wire \mod.flipflop35.q ;
 wire \mod.flipflop36.q ;
 wire \mod.flipflop37.d ;
 wire \mod.flipflop37.q ;
 wire \mod.flipflop38.q ;
 wire \mod.flipflop39.q ;
 wire \mod.flipflop4.q ;
 wire \mod.flipflop40.q ;
 wire \mod.flipflop41.d ;
 wire \mod.flipflop41.q ;
 wire \mod.flipflop42.q ;
 wire \mod.flipflop43.q ;
 wire \mod.flipflop44.q ;
 wire \mod.flipflop45.q ;
 wire \mod.flipflop5.q ;
 wire \mod.flipflop6.q ;
 wire \mod.flipflop8.d ;
 wire \mod.flipflop8.q ;
 wire \mod.flipflop9.d ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;

 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _154_ (.I(\mod.flipflop43.q ),
    .Z(_130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _155_ (.I(_130_),
    .Z(_131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _156_ (.A1(\mod.flipflop11.d ),
    .A2(\mod.flipflop8.q ),
    .Z(_132_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _157_ (.A1(\mod.flipflop33.q ),
    .A2(_131_),
    .A3(_132_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _158_ (.I(_133_),
    .Z(\mod.flipflop8.d ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _159_ (.I(\mod.flipflop40.q ),
    .Z(_134_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _160_ (.A1(\mod.flipflop34.q ),
    .A2(\mod.flipflop35.q ),
    .A3(\mod.flipflop36.q ),
    .A4(\mod.flipflop37.q ),
    .Z(_135_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _161_ (.A1(\mod.flipflop30.q ),
    .A2(\mod.flipflop31.q ),
    .A3(\mod.flipflop32.q ),
    .A4(\mod.flipflop33.q ),
    .ZN(_136_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _162_ (.A1(\mod.flipflop26.q ),
    .A2(\mod.flipflop27.q ),
    .A3(\mod.flipflop28.q ),
    .A4(\mod.flipflop29.q ),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _163_ (.A1(\mod.flipflop38.q ),
    .A2(\mod.flipflop39.q ),
    .A3(\mod.flipflop40.q ),
    .A4(\mod.flipflop41.q ),
    .ZN(_138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _164_ (.A1(_136_),
    .A2(_137_),
    .A3(_138_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _165_ (.A1(\mod.flipflop11.d ),
    .A2(\mod.flipflop8.q ),
    .A3(\mod.flipflop11.q ),
    .A4(\mod.flipflop14.q ),
    .Z(_140_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _166_ (.A1(\mod.flipflop19.q ),
    .A2(\mod.flipflop20.q ),
    .A3(\mod.flipflop22.q ),
    .A4(\mod.flipflop25.q ),
    .ZN(_141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _167_ (.I(\mod.flipflop42.q ),
    .Z(_142_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _168_ (.A1(\mod.flipflop12.q ),
    .A2(\mod.flipflop13.q ),
    .A3(_142_),
    .A4(_130_),
    .ZN(_143_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _169_ (.A1(\mod.flipflop18.q ),
    .A2(\mod.flipflop21.q ),
    .A3(\mod.flipflop23.q ),
    .A4(\mod.flipflop24.q ),
    .ZN(_144_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _170_ (.A1(_141_),
    .A2(_143_),
    .A3(_144_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _171_ (.A1(_135_),
    .A2(_139_),
    .A3(_140_),
    .A4(_145_),
    .ZN(_146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _172_ (.I(_146_),
    .Z(_147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _173_ (.I(_147_),
    .Z(_148_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _174_ (.A1(_134_),
    .A2(_148_),
    .Z(_149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _175_ (.I(_149_),
    .Z(\mod.flipflop41.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _176_ (.A1(\mod.flipflop36.q ),
    .A2(_148_),
    .Z(_150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _177_ (.I(_150_),
    .Z(\mod.flipflop37.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _178_ (.A1(\mod.flipflop33.q ),
    .A2(_148_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _179_ (.I(_151_),
    .Z(\mod.flipflop34.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _180_ (.A1(\mod.flipflop32.q ),
    .A2(_148_),
    .Z(_152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _181_ (.I(_152_),
    .Z(\mod.flipflop33.d ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _182_ (.I(_146_),
    .Z(_153_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _183_ (.A1(\mod.flipflop31.q ),
    .A2(_153_),
    .Z(_000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _184_ (.I(_000_),
    .Z(\mod.flipflop32.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _185_ (.A1(\mod.flipflop28.q ),
    .A2(_153_),
    .Z(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _186_ (.I(_001_),
    .Z(\mod.flipflop29.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _187_ (.A1(\mod.flipflop26.q ),
    .A2(_153_),
    .Z(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _188_ (.I(_002_),
    .Z(\mod.flipflop27.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _189_ (.A1(\mod.flipflop20.q ),
    .A2(_153_),
    .Z(_003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _190_ (.I(_003_),
    .Z(\mod.flipflop21.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _191_ (.A1(\mod.flipflop14.q ),
    .A2(_147_),
    .Z(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _192_ (.I(_004_),
    .Z(\mod.flipflop18.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _193_ (.A1(\mod.flipflop11.q ),
    .A2(_147_),
    .Z(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _194_ (.I(_005_),
    .Z(\mod.flipflop12.d ));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _195_ (.A1(\mod.flipflop8.q ),
    .A2(_147_),
    .Z(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _196_ (.I(_006_),
    .Z(\mod.flipflop9.d ));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _197_ (.A1(\mod.flipflop2.q ),
    .A2(\mod.flipflop3.q ),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _198_ (.A1(\mod.flipflop4.q ),
    .A2(\mod.flipflop5.q ),
    .A3(\mod.flipflop6.q ),
    .A4(\mod.flipflop1.d ),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _199_ (.A1(_007_),
    .A2(_008_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _200_ (.A1(\mod.flipflop44.q ),
    .A2(\mod.flipflop1.q ),
    .A3(\mod.flipflop45.q ),
    .A4(_009_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _201_ (.A1(net15),
    .A2(_010_),
    .Z(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _202_ (.I(_011_),
    .Z(\mod.flipflop2.d ));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _203_ (.I0(net9),
    .I1(net10),
    .I2(net11),
    .I3(net12),
    .S0(\mod.flipflop42.q ),
    .S1(_130_),
    .Z(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _204_ (.I(_012_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _205_ (.I0(net10),
    .I1(net11),
    .I2(net12),
    .I3(net6),
    .S0(\mod.flipflop42.q ),
    .S1(_130_),
    .Z(_014_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _206_ (.I0(net5),
    .I1(net9),
    .I2(net10),
    .I3(net11),
    .S0(\mod.flipflop42.q ),
    .S1(\mod.flipflop43.q ),
    .Z(_015_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _207_ (.A1(_014_),
    .A2(_015_),
    .Z(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _208_ (.I(net8),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _209_ (.I(_017_),
    .Z(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _210_ (.I(net7),
    .Z(_019_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _211_ (.A1(_018_),
    .A2(_019_),
    .Z(_020_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _212_ (.A1(_013_),
    .A2(_016_),
    .A3(_020_),
    .Z(_021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _213_ (.I(_021_),
    .Z(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _214_ (.I(net4),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _215_ (.I(net3),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _216_ (.A1(_023_),
    .A2(_024_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _217_ (.A1(_022_),
    .A2(_025_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _218_ (.I(net2),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _219_ (.A1(_024_),
    .A2(_027_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _220_ (.I(_014_),
    .Z(_029_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _221_ (.A1(_019_),
    .A2(_029_),
    .Z(_030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _222_ (.A1(_019_),
    .A2(_029_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _223_ (.A1(_018_),
    .A2(_012_),
    .Z(_032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _224_ (.I(_015_),
    .Z(_033_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _225_ (.A1(_029_),
    .A2(_033_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _226_ (.A1(_030_),
    .A2(_031_),
    .A3(_032_),
    .B1(_034_),
    .B2(_018_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _227_ (.A1(net4),
    .A2(_028_),
    .B(_035_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _228_ (.A1(_026_),
    .A2(_036_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _229_ (.A1(\mod.flipflop41.q ),
    .A2(_037_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _230_ (.I(_023_),
    .Z(_039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _231_ (.I(_027_),
    .Z(_040_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _232_ (.A1(_039_),
    .A2(_040_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _233_ (.A1(_014_),
    .A2(_033_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _234_ (.I0(_016_),
    .I1(_042_),
    .S(_013_),
    .Z(_043_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _235_ (.A1(_012_),
    .A2(_014_),
    .A3(_033_),
    .Z(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _236_ (.A1(_017_),
    .A2(_044_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _237_ (.A1(_012_),
    .A2(_029_),
    .A3(_033_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _238_ (.A1(_046_),
    .A2(_044_),
    .B(net7),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _239_ (.A1(net8),
    .A2(net7),
    .A3(_043_),
    .B1(_045_),
    .B2(_047_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _240_ (.I(_048_),
    .Z(_049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _241_ (.A1(_023_),
    .A2(net3),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _242_ (.I(_050_),
    .Z(_051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _243_ (.A1(_049_),
    .A2(_051_),
    .B(_022_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _244_ (.A1(_041_),
    .A2(_052_),
    .Z(_053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _245_ (.I(_050_),
    .Z(_054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _246_ (.A1(_049_),
    .A2(_054_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _247_ (.A1(_013_),
    .A2(_016_),
    .A3(_020_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _248_ (.A1(_056_),
    .A2(_025_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _249_ (.I(_057_),
    .Z(_058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _250_ (.I(_035_),
    .Z(_059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _251_ (.I(net2),
    .Z(_060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _252_ (.A1(_023_),
    .A2(net3),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _253_ (.A1(_060_),
    .A2(_061_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _254_ (.A1(_059_),
    .A2(_062_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _255_ (.A1(_055_),
    .A2(_058_),
    .A3(_063_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _256_ (.I(net3),
    .Z(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _257_ (.A1(net4),
    .A2(_027_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _258_ (.A1(_065_),
    .A2(_049_),
    .A3(_066_),
    .Z(_067_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _259_ (.I(_134_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _260_ (.A1(_053_),
    .A2(_064_),
    .A3(_067_),
    .B(_068_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _261_ (.A1(_055_),
    .A2(_057_),
    .A3(_063_),
    .Z(_070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _262_ (.A1(_041_),
    .A2(_052_),
    .B(_067_),
    .ZN(_071_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _263_ (.A1(_134_),
    .A2(_070_),
    .A3(_071_),
    .ZN(_072_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _264_ (.A1(_069_),
    .A2(_072_),
    .Z(_073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _265_ (.A1(_040_),
    .A2(_051_),
    .B(_028_),
    .ZN(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _266_ (.I(_060_),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _267_ (.A1(_075_),
    .A2(_021_),
    .A3(_051_),
    .ZN(_076_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _268_ (.A1(_060_),
    .A2(_025_),
    .ZN(_077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _269_ (.A1(_028_),
    .A2(_077_),
    .ZN(_078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _270_ (.A1(_048_),
    .A2(_062_),
    .B1(_078_),
    .B2(_035_),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _271_ (.A1(_022_),
    .A2(_074_),
    .B(_076_),
    .C(_079_),
    .ZN(_080_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _272_ (.A1(\mod.flipflop39.q ),
    .A2(_080_),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _273_ (.I(_048_),
    .Z(_082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _274_ (.A1(net4),
    .A2(_027_),
    .ZN(_083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _275_ (.A1(_061_),
    .A2(_083_),
    .B1(_077_),
    .B2(_056_),
    .ZN(_084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _276_ (.A1(_082_),
    .A2(_054_),
    .B1(_066_),
    .B2(_059_),
    .C(_084_),
    .ZN(_085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _277_ (.A1(\mod.flipflop35.q ),
    .A2(_085_),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _278_ (.A1(_039_),
    .A2(_075_),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _279_ (.A1(_040_),
    .A2(_061_),
    .B(_035_),
    .ZN(_088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _280_ (.A1(_039_),
    .A2(_060_),
    .ZN(_089_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _281_ (.A1(_039_),
    .A2(_065_),
    .A3(_022_),
    .B(_089_),
    .ZN(_090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _282_ (.A1(_059_),
    .A2(_087_),
    .B(_088_),
    .C(_090_),
    .ZN(_091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _283_ (.A1(_065_),
    .A2(_082_),
    .ZN(_092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _284_ (.A1(\mod.flipflop35.q ),
    .A2(_085_),
    .B1(_091_),
    .B2(_092_),
    .C(\mod.flipflop34.q ),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _285_ (.A1(_024_),
    .A2(_075_),
    .ZN(_094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _286_ (.A1(_075_),
    .A2(_051_),
    .B(_094_),
    .ZN(_095_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _287_ (.A1(_089_),
    .A2(_083_),
    .B(_065_),
    .ZN(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _288_ (.I(_096_),
    .ZN(_097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _289_ (.I0(_095_),
    .I1(_097_),
    .S(_049_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _290_ (.A1(\mod.flipflop36.q ),
    .A2(_058_),
    .A3(_098_),
    .ZN(_099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _291_ (.A1(_086_),
    .A2(_093_),
    .B(_099_),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _292_ (.I(\mod.flipflop37.q ),
    .ZN(_101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _293_ (.A1(_054_),
    .A2(_062_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _294_ (.A1(_040_),
    .A2(_054_),
    .ZN(_103_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _295_ (.A1(_082_),
    .A2(_102_),
    .B(_103_),
    .C(_058_),
    .ZN(_104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _296_ (.A1(_058_),
    .A2(_098_),
    .B(\mod.flipflop36.q ),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _297_ (.A1(_101_),
    .A2(_104_),
    .B(_105_),
    .ZN(_106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _298_ (.A1(_041_),
    .A2(_082_),
    .B1(_092_),
    .B2(_087_),
    .C1(_062_),
    .C2(_059_),
    .ZN(_107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _299_ (.A1(_101_),
    .A2(_104_),
    .ZN(_108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _300_ (.A1(_100_),
    .A2(_106_),
    .B1(_107_),
    .B2(\mod.flipflop38.q ),
    .C(_108_),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _301_ (.A1(_038_),
    .A2(_073_),
    .A3(_081_),
    .A4(_109_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _302_ (.A1(_069_),
    .A2(_072_),
    .A3(_038_),
    .A4(_080_),
    .ZN(_111_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _303_ (.A1(\mod.flipflop38.q ),
    .A2(_107_),
    .Z(_112_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _304_ (.A1(_069_),
    .A2(_072_),
    .A3(_038_),
    .A4(_081_),
    .ZN(_113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _305_ (.A1(_070_),
    .A2(_071_),
    .B(_134_),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _306_ (.A1(_018_),
    .A2(_034_),
    .B1(_043_),
    .B2(_019_),
    .C(_047_),
    .ZN(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _307_ (.I(_115_),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _308_ (.A1(_026_),
    .A2(_036_),
    .B(\mod.flipflop41.q ),
    .ZN(_117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _309_ (.A1(_114_),
    .A2(_038_),
    .B(_116_),
    .C(_117_),
    .ZN(_118_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _310_ (.A1(\mod.flipflop39.q ),
    .A2(_111_),
    .B1(_112_),
    .B2(_113_),
    .C(_118_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _311_ (.A1(_110_),
    .A2(_119_),
    .B(_142_),
    .C(_131_),
    .ZN(_120_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _312_ (.A1(net12),
    .A2(_120_),
    .ZN(_121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _313_ (.I(_121_),
    .Z(\mod.flipflop17.d ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _314_ (.I(_142_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _315_ (.A1(_110_),
    .A2(_119_),
    .B(_122_),
    .C(_131_),
    .ZN(_123_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _316_ (.A1(net11),
    .A2(_123_),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _317_ (.I(_124_),
    .Z(\mod.flipflop16.d ));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _318_ (.I(_131_),
    .ZN(_125_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _319_ (.A1(_110_),
    .A2(_119_),
    .B(_142_),
    .C(_125_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _320_ (.A1(net10),
    .A2(_126_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _321_ (.I(_127_),
    .Z(\mod.flipflop15.d ));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _322_ (.A1(_110_),
    .A2(_119_),
    .B(_122_),
    .C(_125_),
    .ZN(_128_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _323_ (.A1(net9),
    .A2(_128_),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _324_ (.I(_129_),
    .Z(\mod.flipflop10.d ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _325_ (.D(\mod.flipflop37.d ),
    .CLK(net1),
    .Q(\mod.flipflop37.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _326_ (.D(\mod.flipflop35.q ),
    .CLK(net1),
    .Q(\mod.flipflop36.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _327_ (.D(\mod.flipflop34.q ),
    .CLK(net1),
    .Q(\mod.flipflop35.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _328_ (.D(\mod.flipflop34.d ),
    .CLK(net1),
    .Q(\mod.flipflop34.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _329_ (.D(\mod.flipflop33.d ),
    .CLK(net1),
    .Q(\mod.flipflop33.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _330_ (.D(\mod.flipflop32.d ),
    .CLK(net1),
    .Q(\mod.flipflop32.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _331_ (.D(\mod.flipflop30.q ),
    .CLK(net1),
    .Q(\mod.flipflop31.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _332_ (.D(\mod.flipflop29.q ),
    .CLK(net1),
    .Q(\mod.flipflop30.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _333_ (.D(\mod.flipflop29.d ),
    .CLK(net1),
    .Q(\mod.flipflop29.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _334_ (.D(\mod.flipflop27.q ),
    .CLK(net1),
    .Q(\mod.flipflop28.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _335_ (.D(\mod.flipflop27.d ),
    .CLK(net1),
    .Q(\mod.flipflop27.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _336_ (.D(\mod.flipflop25.q ),
    .CLK(net1),
    .Q(\mod.flipflop26.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _337_ (.D(\mod.flipflop24.q ),
    .CLK(net1),
    .Q(\mod.flipflop25.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _338_ (.D(\mod.flipflop23.q ),
    .CLK(net1),
    .Q(\mod.flipflop24.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _339_ (.D(\mod.flipflop22.q ),
    .CLK(net1),
    .Q(\mod.flipflop23.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _340_ (.D(\mod.flipflop21.q ),
    .CLK(net1),
    .Q(\mod.flipflop22.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _341_ (.D(\mod.flipflop21.d ),
    .CLK(net1),
    .Q(\mod.flipflop21.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _342_ (.D(\mod.flipflop19.q ),
    .CLK(net1),
    .Q(\mod.flipflop20.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _343_ (.D(\mod.flipflop18.q ),
    .CLK(net1),
    .Q(\mod.flipflop19.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _344_ (.D(\mod.flipflop18.d ),
    .CLK(net1),
    .Q(\mod.flipflop18.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _345_ (.D(\mod.flipflop13.q ),
    .CLK(net1),
    .Q(\mod.flipflop14.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _346_ (.D(\mod.flipflop12.q ),
    .CLK(net1),
    .Q(\mod.flipflop13.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _347_ (.D(\mod.flipflop12.d ),
    .CLK(net1),
    .Q(\mod.flipflop12.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _348_ (.D(\mod.flipflop11.d ),
    .CLK(net1),
    .Q(\mod.flipflop11.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _349_ (.D(\mod.flipflop9.d ),
    .CLK(net1),
    .Q(\mod.flipflop11.d ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _350_ (.D(\mod.flipflop8.d ),
    .CLK(net1),
    .Q(\mod.flipflop8.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _351_ (.D(\mod.flipflop6.q ),
    .CLK(net1),
    .Q(\mod.flipflop1.d ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _352_ (.D(\mod.flipflop5.q ),
    .CLK(net1),
    .Q(\mod.flipflop6.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _353_ (.D(\mod.flipflop4.q ),
    .CLK(net1),
    .Q(\mod.flipflop5.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _354_ (.D(\mod.flipflop3.q ),
    .CLK(net1),
    .Q(\mod.flipflop4.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _355_ (.D(\mod.flipflop2.q ),
    .CLK(net1),
    .Q(\mod.flipflop3.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _356_ (.D(\mod.flipflop2.d ),
    .CLK(net1),
    .Q(\mod.flipflop2.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _357_ (.D(\mod.flipflop17.d ),
    .CLK(net15),
    .Q(net12));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _358_ (.D(\mod.flipflop16.d ),
    .CLK(net15),
    .Q(net11));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _359_ (.D(\mod.flipflop15.d ),
    .CLK(net15),
    .Q(net10));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _360_ (.D(\mod.flipflop10.d ),
    .CLK(net15),
    .Q(net9));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _361_ (.D(\mod.flipflop45.q ),
    .CLK(net1),
    .Q(net15));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _362_ (.D(\mod.flipflop44.q ),
    .CLK(net1),
    .Q(\mod.flipflop45.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _363_ (.D(\mod.flipflop1.q ),
    .CLK(net1),
    .Q(\mod.flipflop44.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _364_ (.D(\mod.flipflop1.d ),
    .CLK(net1),
    .Q(\mod.flipflop1.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _365_ (.D(\mod.flipflop42.q ),
    .CLK(net1),
    .Q(\mod.flipflop43.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _366_ (.D(\mod.flipflop41.q ),
    .CLK(net1),
    .Q(\mod.flipflop42.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _367_ (.D(\mod.flipflop41.d ),
    .CLK(net1),
    .Q(\mod.flipflop41.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _368_ (.D(\mod.flipflop39.q ),
    .CLK(net1),
    .Q(\mod.flipflop40.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _369_ (.D(\mod.flipflop38.q ),
    .CLK(net1),
    .Q(\mod.flipflop39.q ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _370_ (.D(\mod.flipflop37.q ),
    .CLK(net1),
    .Q(\mod.flipflop38.q ));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_17 (.ZN(net17));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_18 (.ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_19 (.ZN(net19));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_20 (.ZN(net20));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_21 (.ZN(net21));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_22 (.ZN(net22));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_23 (.ZN(net23));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_24 (.ZN(net24));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_25 (.ZN(net25));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_26 (.ZN(net26));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_27 (.ZN(net27));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_28 (.ZN(net28));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_29 (.ZN(net29));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_30 (.ZN(net30));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_31 (.ZN(net31));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_32 (.ZN(net32));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_33 (.ZN(net33));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_34 (.ZN(net34));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_35 (.ZN(net35));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_36 (.ZN(net36));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_37 (.ZN(net37));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_38 (.ZN(net38));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_39 (.ZN(net39));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_40 (.ZN(net40));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_41 (.ZN(net41));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_42 (.ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_43 (.ZN(net43));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_44 (.ZN(net44));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_45 (.ZN(net45));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_46 (.ZN(net46));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_47 (.ZN(net47));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_48 (.ZN(net48));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_49 (.ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_50 (.ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_51 (.ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_52 (.ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__186__I (.I(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _440_ (.I(net6),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _441_ (.I(net5),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 input1 (.I(io_in[12]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(io_in[13]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(io_in[14]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(io_in[15]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(io_in[16]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(io_in[17]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(io_in[18]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[19]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output9 (.I(net9),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output10 (.I(net10),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output11 (.I(net11),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output12 (.I(net12),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output13 (.I(net13),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output14 (.I(net14),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 output15 (.I(net15),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__tiel tiny_user_project_16 (.ZN(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__190__I (.I(_003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__192__I (.I(_004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__194__I (.I(_005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__196__I (.I(_006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__A1 (.I(_007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__199__A2 (.I(_008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__202__I (.I(_011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__A1 (.I(_012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__A1 (.I(_012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__A2 (.I(_012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__204__I (.I(_012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A1 (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__S (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__A1 (.I(_013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__A2 (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__A1 (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__220__I (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__207__A1 (.I(_014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__224__I (.I(_015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__207__A2 (.I(_015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A2 (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__I0 (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__A2 (.I(_016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__A1 (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__209__I (.I(_017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__A1 (.I(_018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__B2 (.I(_018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__223__A1 (.I(_018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__A1 (.I(_018_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__B2 (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__A1 (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__221__A1 (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__211__A2 (.I(_019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__247__A3 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__212__A3 (.I(_020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__A3 (.I(_022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__A1 (.I(_022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__B (.I(_022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__A1 (.I(_022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__A1 (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__A1 (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__230__I (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__A1 (.I(_023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__A1 (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__A1 (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__216__A2 (.I(_024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__A2 (.I(_025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__A2 (.I(_025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__217__A2 (.I(_025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__A1 (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__A1 (.I(_026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__274__A2 (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__A2 (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__231__I (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__219__A2 (.I(_027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__A1 (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__B (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__A2 (.I(_028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__A2 (.I(_029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__225__A1 (.I(_029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__222__A2 (.I(_029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__221__A2 (.I(_029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__A1 (.I(_030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__A2 (.I(_031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__A3 (.I(_032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__237__A3 (.I(_033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__235__A3 (.I(_033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__233__A2 (.I(_033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__225__A2 (.I(_033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__A2 (.I(_034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__226__B1 (.I(_034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__B (.I(_035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__B2 (.I(_035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__250__I (.I(_035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__B (.I(_035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__228__A2 (.I(_036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__A2 (.I(_037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__A2 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A3 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A3 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__A1 (.I(_038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__A1 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__A1 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A1 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__A1 (.I(_039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__A1 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__A1 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__A1 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__232__A2 (.I(_040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__A1 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A1 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__244__A1 (.I(_041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__234__I1 (.I(_042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__B1 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__A3 (.I(_043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__A2 (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__236__A2 (.I(_044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__A1 (.I(_046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__306__C (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__B2 (.I(_047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__S (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A2 (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__A1 (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__A1 (.I(_049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__245__I (.I(_050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__242__I (.I(_050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__A2 (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__A3 (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__265__A2 (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__243__A2 (.I(_051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__A2 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__244__A2 (.I(_052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A1 (.I(_053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__294__A2 (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A1 (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__A2 (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__246__A2 (.I(_054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__A1 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__A1 (.I(_055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__B2 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__248__A1 (.I(_056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__A2 (.I(_057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__249__I (.I(_057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A1 (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__C (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A2 (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__A2 (.I(_058_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__C2 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__B2 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__A1 (.I(_059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__280__A2 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__268__A1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__266__I (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__A1 (.I(_060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__279__A2 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A1 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__253__A2 (.I(_061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__C1 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__293__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__270__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__254__A2 (.I(_062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__261__A3 (.I(_063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__255__A3 (.I(_063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A2 (.I(_064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__B (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__A1 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__A2 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A1 (.I(_065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__B1 (.I(_066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__258__A3 (.I(_066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__262__B (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__A3 (.I(_067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__260__B (.I(_068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__A1 (.I(_069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__A2 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__A2 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__A3 (.I(_071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A2 (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A2 (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__264__A2 (.I(_072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__A2 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__A2 (.I(_074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__A1 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__285__A2 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__278__A2 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__267__A1 (.I(_075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__271__B (.I(_076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__B1 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__269__A2 (.I(_077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__302__A4 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A2 (.I(_080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__304__A4 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__A3 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__A2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__283__A2 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__A1 (.I(_082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A2 (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__275__A2 (.I(_083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__276__C (.I(_084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A2 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__A2 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__B2 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__A2 (.I(_087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__282__B (.I(_088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__287__A1 (.I(_089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__281__B (.I(_089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__B1 (.I(_091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__298__B1 (.I(_092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__B2 (.I(_092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__291__A2 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__286__B (.I(_094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__I0 (.I(_095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__289__I1 (.I(_097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__A2 (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A3 (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__A1 (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A1 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A1 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__295__A2 (.I(_102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__299__A2 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__A2 (.I(_104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__297__B (.I(_105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A2 (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__B1 (.I(_107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__C (.I(_108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__301__A4 (.I(_109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__B1 (.I(_112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__A1 (.I(_114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__309__B (.I(_116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__A2 (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__A2 (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__A2 (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__A2 (.I(_119_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__A2 (.I(_120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__313__I (.I(_121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__B (.I(_122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__B (.I(_122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A2 (.I(_123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__322__C (.I(_125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__C (.I(_125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__321__I (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__324__I (.I(_129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__S1 (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__S1 (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__A4 (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__155__I (.I(_130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__318__I (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__315__C (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__C (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__A2 (.I(_131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__305__B (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__263__A1 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__259__I (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__A1 (.I(_134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__A1 (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__A1 (.I(_136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__164__A2 (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__170__A1 (.I(_141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__319__B (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__314__I (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__311__B (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__A3 (.I(_142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__171__A4 (.I(_145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__182__I (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__172__I (.I(_146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__A2 (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__193__A2 (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__191__A2 (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__173__I (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__A2 (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__A2 (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__A2 (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__174__A2 (.I(_148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__175__I (.I(_149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__177__I (.I(_150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__179__I (.I(_151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__181__I (.I(_152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__A2 (.I(_153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__A2 (.I(_153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__A2 (.I(_153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__A2 (.I(_153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[16]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[17]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[18]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[19]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__D (.I(\mod.flipflop1.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__198__A4 (.I(\mod.flipflop1.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__D (.I(\mod.flipflop1.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__A2 (.I(\mod.flipflop1.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__D (.I(\mod.flipflop10.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__D (.I(\mod.flipflop11.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__A1 (.I(\mod.flipflop11.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__A1 (.I(\mod.flipflop11.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__193__A1 (.I(\mod.flipflop11.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__A3 (.I(\mod.flipflop11.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__D (.I(\mod.flipflop12.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__D (.I(\mod.flipflop12.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__A1 (.I(\mod.flipflop12.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__D (.I(\mod.flipflop13.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__168__A2 (.I(\mod.flipflop13.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__191__A1 (.I(\mod.flipflop14.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__A4 (.I(\mod.flipflop14.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__D (.I(\mod.flipflop16.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__D (.I(\mod.flipflop17.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__D (.I(\mod.flipflop18.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__A1 (.I(\mod.flipflop18.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__D (.I(\mod.flipflop19.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__166__A1 (.I(\mod.flipflop19.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__D (.I(\mod.flipflop2.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__D (.I(\mod.flipflop2.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__A1 (.I(\mod.flipflop2.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__189__A1 (.I(\mod.flipflop20.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__166__A2 (.I(\mod.flipflop20.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__D (.I(\mod.flipflop21.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__D (.I(\mod.flipflop21.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__A2 (.I(\mod.flipflop21.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__D (.I(\mod.flipflop22.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__166__A3 (.I(\mod.flipflop22.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__D (.I(\mod.flipflop23.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__A3 (.I(\mod.flipflop23.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__D (.I(\mod.flipflop24.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__169__A4 (.I(\mod.flipflop24.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__D (.I(\mod.flipflop25.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__166__A4 (.I(\mod.flipflop25.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__187__A1 (.I(\mod.flipflop26.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__A1 (.I(\mod.flipflop26.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__D (.I(\mod.flipflop27.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__185__A1 (.I(\mod.flipflop28.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__162__A3 (.I(\mod.flipflop28.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__D (.I(\mod.flipflop29.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__D (.I(\mod.flipflop3.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__197__A2 (.I(\mod.flipflop3.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__D (.I(\mod.flipflop30.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__A1 (.I(\mod.flipflop30.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__183__A1 (.I(\mod.flipflop31.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__A2 (.I(\mod.flipflop31.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__D (.I(\mod.flipflop32.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__180__A1 (.I(\mod.flipflop32.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__A3 (.I(\mod.flipflop32.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__D (.I(\mod.flipflop33.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__178__A1 (.I(\mod.flipflop33.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__161__A4 (.I(\mod.flipflop33.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__157__A1 (.I(\mod.flipflop33.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__D (.I(\mod.flipflop34.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__D (.I(\mod.flipflop34.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__C (.I(\mod.flipflop34.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__A1 (.I(\mod.flipflop34.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__D (.I(\mod.flipflop35.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__284__A1 (.I(\mod.flipflop35.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__277__A1 (.I(\mod.flipflop35.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__A2 (.I(\mod.flipflop35.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__296__B (.I(\mod.flipflop36.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__290__A1 (.I(\mod.flipflop36.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__176__A1 (.I(\mod.flipflop36.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__A3 (.I(\mod.flipflop36.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__D (.I(\mod.flipflop37.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__D (.I(\mod.flipflop37.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__292__I (.I(\mod.flipflop37.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__160__A4 (.I(\mod.flipflop37.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__D (.I(\mod.flipflop38.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__303__A1 (.I(\mod.flipflop38.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__300__B2 (.I(\mod.flipflop38.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__A1 (.I(\mod.flipflop38.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__D (.I(\mod.flipflop39.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__310__A1 (.I(\mod.flipflop39.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__272__A1 (.I(\mod.flipflop39.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__A2 (.I(\mod.flipflop39.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__D (.I(\mod.flipflop4.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__198__A1 (.I(\mod.flipflop4.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__A3 (.I(\mod.flipflop40.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__159__I (.I(\mod.flipflop40.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__D (.I(\mod.flipflop41.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__D (.I(\mod.flipflop41.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__308__B (.I(\mod.flipflop41.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__229__A1 (.I(\mod.flipflop41.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__163__A4 (.I(\mod.flipflop41.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__D (.I(\mod.flipflop42.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__S0 (.I(\mod.flipflop42.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__S0 (.I(\mod.flipflop42.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__S0 (.I(\mod.flipflop42.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__167__I (.I(\mod.flipflop42.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__S1 (.I(\mod.flipflop43.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__154__I (.I(\mod.flipflop43.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__D (.I(\mod.flipflop44.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__A1 (.I(\mod.flipflop44.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__D (.I(\mod.flipflop45.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__200__A3 (.I(\mod.flipflop45.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__D (.I(\mod.flipflop5.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__198__A2 (.I(\mod.flipflop5.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__D (.I(\mod.flipflop8.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__195__A1 (.I(\mod.flipflop8.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__165__A2 (.I(\mod.flipflop8.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__156__A2 (.I(\mod.flipflop8.q ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__D (.I(\mod.flipflop9.d ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__370__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__369__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__368__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__367__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__366__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__365__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__364__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__363__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__362__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__361__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__356__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__355__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__354__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__353__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__352__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__351__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__350__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__349__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__348__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__347__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__346__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__345__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__344__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__343__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__342__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__341__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__340__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__339__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__338__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__337__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__336__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__335__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__334__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__333__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__332__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__331__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__330__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__329__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__328__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__327__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__326__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__325__CLK (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__251__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__218__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__256__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__252__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__241__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__215__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__274__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__257__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__227__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__214__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I0 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__440__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__I3 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__239__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__238__B (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__210__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output9_I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__323__A1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I1 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I0 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output10_I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__320__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__I0 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__316__A1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__206__I3 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__I1 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__312__A1 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__205__I2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__203__I3 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__360__CLK (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__359__CLK (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__358__CLK (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__357__CLK (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__201__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_5_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_5_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_6_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_7_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_7_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_8_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_8_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_9_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_9_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_10_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_11_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_11_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_12_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_13_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_13_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_14_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_15_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_15_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_16_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_17_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_17_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_18_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_18_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_19_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_19_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_20_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_21_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_21_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_22_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_26_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_27_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_27_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_28_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_29_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_29_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_30_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_30_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_31_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_31_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_32_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_32_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_33_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_33_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_34_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_35_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_35_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_36_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_37_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_38_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_39_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_40_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_40_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_41_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_41_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_419 ();
 assign io_oeb[0] = net52;
 assign io_oeb[10] = net62;
 assign io_oeb[11] = net63;
 assign io_oeb[12] = net64;
 assign io_oeb[13] = net65;
 assign io_oeb[14] = net66;
 assign io_oeb[15] = net67;
 assign io_oeb[16] = net68;
 assign io_oeb[17] = net69;
 assign io_oeb[18] = net70;
 assign io_oeb[19] = net71;
 assign io_oeb[1] = net53;
 assign io_oeb[20] = net72;
 assign io_oeb[21] = net73;
 assign io_oeb[22] = net74;
 assign io_oeb[23] = net75;
 assign io_oeb[24] = net76;
 assign io_oeb[25] = net77;
 assign io_oeb[26] = net78;
 assign io_oeb[27] = net79;
 assign io_oeb[28] = net80;
 assign io_oeb[29] = net81;
 assign io_oeb[2] = net54;
 assign io_oeb[30] = net82;
 assign io_oeb[31] = net83;
 assign io_oeb[32] = net84;
 assign io_oeb[33] = net16;
 assign io_oeb[34] = net17;
 assign io_oeb[35] = net18;
 assign io_oeb[36] = net19;
 assign io_oeb[37] = net20;
 assign io_oeb[3] = net55;
 assign io_oeb[4] = net56;
 assign io_oeb[5] = net57;
 assign io_oeb[6] = net58;
 assign io_oeb[7] = net59;
 assign io_oeb[8] = net60;
 assign io_oeb[9] = net61;
 assign io_out[0] = net21;
 assign io_out[10] = net31;
 assign io_out[11] = net32;
 assign io_out[12] = net33;
 assign io_out[13] = net34;
 assign io_out[14] = net35;
 assign io_out[15] = net36;
 assign io_out[16] = net37;
 assign io_out[17] = net38;
 assign io_out[18] = net39;
 assign io_out[19] = net40;
 assign io_out[1] = net22;
 assign io_out[26] = net41;
 assign io_out[28] = net42;
 assign io_out[29] = net43;
 assign io_out[2] = net23;
 assign io_out[30] = net44;
 assign io_out[31] = net45;
 assign io_out[32] = net46;
 assign io_out[33] = net47;
 assign io_out[34] = net48;
 assign io_out[35] = net49;
 assign io_out[36] = net50;
 assign io_out[37] = net51;
 assign io_out[3] = net24;
 assign io_out[4] = net25;
 assign io_out[5] = net26;
 assign io_out[6] = net27;
 assign io_out[7] = net28;
 assign io_out[8] = net29;
 assign io_out[9] = net30;
endmodule

