* NGSPICE file created from tiny_user_project.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

.subckt tiny_user_project io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vccd1 vssd1
XFILLER_54_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_294_ _040_ _054_ _103_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_363_ mod.flipflop1.q net1 mod.flipflop44.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__249__I _057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__159__I mod.flipflop40.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_346_ mod.flipflop12.q net1 mod.flipflop13.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_277_ mod.flipflop35.q _085_ _086_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_200_ mod.flipflop44.q mod.flipflop1.q mod.flipflop45.q _009_ _010_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__180__A2 _148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__235__A3 _033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_329_ mod.flipflop33.d net1 mod.flipflop33.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__226__A3 _032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__234__I0 _016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__351__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__172__I _146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__167__I mod.flipflop42.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_304 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__283__A1 _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__274__A1 net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_362_ mod.flipflop44.q net1 mod.flipflop45.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_293_ _054_ _062_ _102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__265__A1 _040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__247__A1 _013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_276_ _082_ _054_ _066_ _059_ _084_ _085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__175__I _149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_345_ mod.flipflop13.q net1 mod.flipflop14.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__238__A1 _046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__229__A1 mod.flipflop41.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_328_ mod.flipflop34.d net1 mod.flipflop34.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_259_ _134_ _068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__234__I1 _042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__162__A3 mod.flipflop28.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output12_I net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__310__B1 _112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__206__S0 mod.flipflop42.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_338 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__341__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput10 net10 io_out[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__364__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__289__S _049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input3_I io_in[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__283__A2 _082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_146 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_135 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__274__A2 _027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_361_ mod.flipflop45.q net1 net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_292_ mod.flipflop37.q _101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__265__A2 _051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__247__A2 _016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__183__A1 mod.flipflop31.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_344_ mod.flipflop18.d net1 mod.flipflop18.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_275_ _061_ _083_ _077_ _056_ _084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__238__A2 _044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__315__B _122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__174__A1 _134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__229__A2 _037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__165__A1 mod.flipflop11.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__186__I _001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_327_ mod.flipflop34.q net1 mod.flipflop35.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__171__A4 _145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_258_ _065_ _049_ _066_ _067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_189_ mod.flipflop20.q _153_ _003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__156__A1 mod.flipflop11.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__310__A1 mod.flipflop39.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__301__A1 _038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__206__S1 mod.flipflop43.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_306 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput11 net11 io_out[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput9 net9 io_out[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__194__I _005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_169 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_11_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_291_ _086_ _093_ _099_ _100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_360_ mod.flipflop10.d net15 net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__331__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__354__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__247__A3 _020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__183__A2 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_343_ mod.flipflop18.q net1 mod.flipflop19.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_274_ net4 _027_ _083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__315__C _131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__174__A2 _148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__165__A2 mod.flipflop8.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__292__I mod.flipflop37.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_326_ mod.flipflop35.q net1 mod.flipflop36.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_188_ _002_ mod.flipflop27.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__156__A2 mod.flipflop8.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_257_ net4 _027_ _066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_309_ _114_ _038_ _116_ _117_ _118_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_42_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__301__A2 _073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__295__A1 _082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__286__A1 _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput12 net12 io_out[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__277__A1 mod.flipflop35.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__201__A1 net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__268__A1 _060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_290_ mod.flipflop36.q _058_ _098_ _099_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_342_ mod.flipflop19.q net1 mod.flipflop20.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_273_ _048_ _082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__165__A3 mod.flipflop11.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_325_ mod.flipflop37.d net1 mod.flipflop37.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_14_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_187_ mod.flipflop26.q _153_ _002_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_256_ net3 _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__344__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__367__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_308_ _026_ _036_ mod.flipflop41.q _117_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_239_ net8 net7 _043_ _045_ _047_ _048_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__301__A3 _081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__298__C1 _062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output10_I net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_308 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__295__A2 _102_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_168 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__286__A2 _051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput13 net13 io_out[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__277__A2 _085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_138 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__268__A2 _025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__195__A1 mod.flipflop8.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__260__B _068_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_341_ mod.flipflop21.d net1 mod.flipflop21.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__168__A1 mod.flipflop12.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_272_ mod.flipflop39.q _080_ _081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_49_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__331__D mod.flipflop30.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__165__A4 mod.flipflop14.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__322__A1 _110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_324_ _129_ mod.flipflop10.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_255_ _055_ _058_ _063_ _064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_43_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_186_ _001_ mod.flipflop29.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__326__D mod.flipflop35.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__304__A1 _069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_238_ _046_ _044_ net7 _047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_307_ _115_ _116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_169_ mod.flipflop18.q mod.flipflop21.q mod.flipflop23.q mod.flipflop24.q _144_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__301__A4 _109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__298__C2 _059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__298__B1 _092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__334__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__357__CLK net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput14 net14 io_out[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_44_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_0 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__195__A2 _147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__329__D mod.flipflop33.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_271_ _022_ _074_ _076_ _079_ _080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_340_ mod.flipflop21.q net1 mod.flipflop22.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__168__A2 mod.flipflop13.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__271__B _076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__322__A2 _119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_254_ _059_ _062_ _063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_185_ mod.flipflop28.q _153_ _001_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_13_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_323_ net9 _128_ _129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__342__D mod.flipflop19.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__304__A2 _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_306_ _018_ _034_ _043_ _019_ _047_ _115_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_34_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_237_ _012_ _029_ _033_ _046_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_168_ mod.flipflop12.q mod.flipflop13.q _142_ _130_ _143_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__298__A1 _041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__298__B2 _087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__222__A1 _019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__337__D mod.flipflop24.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput15 net15 io_out[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_35_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__350__D mod.flipflop8.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__347__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__345__D mod.flipflop13.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_270_ _048_ _062_ _078_ _035_ _079_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_41_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__168__A3 _142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_290 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_322_ _110_ _119_ _122_ _125_ _128_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_184_ _000_ mod.flipflop32.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_253_ _060_ _061_ _062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__282__B _088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__304__A3 _038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_305_ _070_ _071_ _134_ _114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_236_ _017_ _044_ _045_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__298__A2 _082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_167_ mod.flipflop42.q _142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__222__A2 _029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__353__D mod.flipflop4.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_219_ _024_ _027_ _028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__348__D mod.flipflop11.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__198__A1 mod.flipflop4.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__189__A1 mod.flipflop20.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__361__D mod.flipflop45.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__214__I net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__168__A4 _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__316__A1 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__356__D mod.flipflop2.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__209__I _017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_291 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_252_ _023_ net3 _061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_321_ _127_ mod.flipflop15.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_183_ mod.flipflop31.q _153_ _000_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_49_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__337__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__304__A4 _081_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_304_ _069_ _072_ _038_ _081_ _113_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_10_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_235_ _012_ _014_ _033_ _044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
X_166_ mod.flipflop19.q mod.flipflop20.q mod.flipflop22.q mod.flipflop25.q _141_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_41_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_158 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_218_ net2 _027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__364__D mod.flipflop1.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__203__I0 net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__198__A2 mod.flipflop5.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__189__A2 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__370__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output9_I net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__230__I _023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__270__B2 _035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__261__A1 _055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__296__B mod.flipflop36.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__316__A2 _123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__252__A1 _023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__243__A1 _049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_320_ net10 _126_ _127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_182_ _146_ _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_251_ net2 _060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_6_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__225__A1 _029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__367__D mod.flipflop41.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__216__A1 _023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_234_ _016_ _042_ _013_ _043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_303_ mod.flipflop38.q _107_ _112_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
X_165_ mod.flipflop11.d mod.flipflop8.q mod.flipflop11.q mod.flipflop14.q _140_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_40_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__207__A1 _014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_126 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__327__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_217_ _022_ _025_ _026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__203__I1 net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_102 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_21_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__318__I _131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__270__A2 _062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__261__A2 _057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__252__A2 net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__360__CLK net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__243__A2 _051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_181_ _152_ mod.flipflop33.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_250_ _035_ _059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__170__A1 _141_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__225__A2 _033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__161__A1 mod.flipflop30.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_302_ _069_ _072_ _038_ _080_ _111_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__216__A2 _024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_233_ _014_ _033_ _042_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_164_ _136_ _137_ _138_ _139_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_49_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__207__A2 _015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_216_ _023_ _024_ _025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__203__I2 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__198__A4 mod.flipflop1.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__154__I mod.flipflop43.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__319__A1 _110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__261__A3 _063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_272 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_294 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_180_ mod.flipflop32.q _148_ _152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_22_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__161__A2 mod.flipflop31.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_301_ _038_ _073_ _081_ _109_ _110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and4_1
X_232_ _039_ _040_ _041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_163_ mod.flipflop38.q mod.flipflop39.q mod.flipflop40.q mod.flipflop41.q _138_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_40_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__350__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__206__I0 net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_215_ net3 _024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__203__I3 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_20_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__440__I net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input8_I io_in[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__282__A1 _059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__264__A1 _069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__319__A2 _119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_421 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_410 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__255__A1 _055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__246__A1 _049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__237__A1 _012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__228__A1 _026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_262 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_284 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__219__A1 _024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__161__A3 mod.flipflop32.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_162_ mod.flipflop26.q mod.flipflop27.q mod.flipflop28.q mod.flipflop29.q _137_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_300_ _100_ _106_ _107_ mod.flipflop38.q _108_ _109_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_10_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_231_ _027_ _040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_118 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__300__B1 _107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 io_in[12] net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_45_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__206__I1 net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__205__S0 mod.flipflop42.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_214_ net4 _023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__173__I _147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__340__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__291__A2 _093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__282__A2 _087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__363__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__264__A2 _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_400 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_422 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__255__A2 _058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__191__A1 mod.flipflop14.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__246__A2 _054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__181__I _152_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__237__A2 _029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__305__B _134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_241 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__228__A2 _036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_296 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__266__I _060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__164__A1 _136_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__219__A2 _027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__161__A4 mod.flipflop33.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_161_ mod.flipflop30.q mod.flipflop31.q mod.flipflop32.q mod.flipflop33.q _136_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_230_ _023_ _039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_359_ mod.flipflop15.d net15 net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_46_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__300__A1 _100_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__300__B2 mod.flipflop38.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 io_in[13] net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__206__I2 net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__205__S1 _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_213_ _021_ _022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_106 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__276__B1 _066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_11_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__308__B mod.flipflop41.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__179__I _151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_401 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__255__A3 _063_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__330__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__191__A2 _147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__237__A3 _033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__353__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_220 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_231 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_253 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__164__A2 _137_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__192__I _004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_160_ mod.flipflop34.q mod.flipflop35.q mod.flipflop36.q mod.flipflop37.q _135_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_49_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_358_ mod.flipflop16.d net15 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_18_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_289_ _095_ _097_ _049_ _098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_39_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput3 io_in[14] net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__206__I3 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output15_I net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_212_ _013_ _016_ _020_ _021_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_30_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__294__A1 _040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_178 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__285__A1 _024_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__276__B2 _059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__276__A1 _082_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__200__A1 mod.flipflop44.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__267__A1 _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__258__A1 _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_251 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_402 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__319__B _142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_221 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_232 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_276 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_287 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_298 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__343__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_357_ mod.flipflop17.d net15 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_288_ _096_ _097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[15] net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__366__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_211_ _018_ _019_ _020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_42_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__294__A2 _054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__285__A2 _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__276__A2 _054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__200__A2 mod.flipflop1.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__258__A2 _049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__185__A1 mod.flipflop28.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__319__C _125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__176__A1 mod.flipflop36.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_200 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_233 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_255 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_266 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_288 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__312__A1 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__303__A1 mod.flipflop38.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_356_ mod.flipflop2.d net1 mod.flipflop2.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_287_ _089_ _083_ _065_ _096_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput5 io_in[16] net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_80 io_oeb[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_210_ net7 _019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_339_ mod.flipflop22.q net1 mod.flipflop23.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__333__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_46_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__200__A3 mod.flipflop45.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__356__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__267__A3 _051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__258__A3 _066_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__185__A2 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_415 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_404 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__176__A2 _148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_201 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_223 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_256 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_267 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_359 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_441_ net5 net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__312__A2 _120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__303__A2 _107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_286_ _075_ _051_ _094_ _095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_355_ mod.flipflop2.q net1 mod.flipflop3.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__297__A1 _101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_70 io_oeb[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput6 io_in[17] net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_81 io_oeb[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_24_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_156 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__327__D mod.flipflop34.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__221__A1 _019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__212__A1 _013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__279__A1 _040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_338_ mod.flipflop23.q net1 mod.flipflop24.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_90 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_269_ _028_ _077_ _078_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output13_I net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__340__D mod.flipflop21.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_7_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__335__D mod.flipflop27.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__346__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_213 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_235 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input4_I io_in[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_268 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__369__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__306__B1 _043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_440_ net6 net13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_13_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_354_ mod.flipflop3.q net1 mod.flipflop4.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_285_ _024_ _075_ _094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__297__A2 _104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xtiny_user_project_71 io_oeb[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xinput7 io_in[18] net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_82 io_oeb[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_60 io_oeb[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__221__A2 _029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__343__D mod.flipflop18.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__212__A2 _016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__279__A2 _061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_91 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_337_ mod.flipflop24.q net1 mod.flipflop25.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_268_ _060_ _025_ _077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_199_ _007_ _008_ _009_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__338__D mod.flipflop23.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__197__A1 mod.flipflop2.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_263 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_274 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_406 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__204__I _012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__315__A1 _110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_203 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_225 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_236 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__346__D mod.flipflop12.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__306__A1 _018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__306__B2 _019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_370_ mod.flipflop37.q net1 mod.flipflop38.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_5_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__336__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_284_ mod.flipflop35.q _085_ _091_ _092_ mod.flipflop34.q _093_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_41_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_353_ mod.flipflop4.q net1 mod.flipflop5.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__359__CLK net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput8 io_in[19] net8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xtiny_user_project_72 io_oeb[20] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_61 io_oeb[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_50 io_out[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_83 io_oeb[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_136 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__212__A3 _020_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_336_ mod.flipflop25.q net1 mod.flipflop26.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_267_ _075_ _021_ _051_ _076_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_198_ mod.flipflop4.q mod.flipflop5.q mod.flipflop6.q mod.flipflop1.d _008_ vccd1
+ vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_32_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__354__D mod.flipflop3.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__197__A2 mod.flipflop3.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_275 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_319_ _110_ _119_ _142_ _125_ _126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__349__D mod.flipflop9.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_407 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__220__I _014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__286__B _094_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__260__A1 _053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__315__A2 _119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_248 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__215__I net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__362__D mod.flipflop44.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__306__A2 _034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_134 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__233__A1 _014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_112 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__357__D mod.flipflop17.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_283_ _065_ _082_ _092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_352_ mod.flipflop5.q net1 mod.flipflop6.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xtiny_user_project_51 io_out[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_84 io_oeb[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_62 io_oeb[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_40 io_out[19] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_73 io_oeb[21] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_148 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_82 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_71 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_197_ mod.flipflop2.q mod.flipflop3.q _007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_335_ mod.flipflop27.d net1 mod.flipflop27.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__326__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_266_ _060_ _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__313__I _121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_295 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__370__D mod.flipflop37.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__349__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_249_ _057_ _058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_318_ _131_ _125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_35_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__365__D mod.flipflop42.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__218__I net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output11_I net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__260__A2 _064_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_205 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__321__I _127_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_216 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_227 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_249 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__231__I _027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__297__B _105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__233__A2 _033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I io_in[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_124 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__160__A1 mod.flipflop34.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_351_ mod.flipflop6.q net1 mod.flipflop1.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_26_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_282_ _059_ _087_ _088_ _090_ _091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_5_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_41 io_out[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_63 io_oeb[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_52 io_oeb[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_74 io_oeb[22] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_30 io_out[9] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__368__D mod.flipflop39.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_334_ mod.flipflop27.q net1 mod.flipflop28.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_83 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_196_ _006_ mod.flipflop9.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_265_ _040_ _051_ _028_ _074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_317_ _124_ mod.flipflop16.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_248_ _056_ _025_ _057_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__324__I _129_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_179_ _151_ mod.flipflop34.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_47_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_214 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__339__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__309__A1 _114_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__260__A3 _067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_217 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_228 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__160__A2 mod.flipflop35.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__242__I _050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_350_ mod.flipflop8.d net1 mod.flipflop8.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_281_ _039_ _065_ _022_ _089_ _090_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_5_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_31 io_out[10] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_20 io_oeb[37] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_53 io_oeb[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_64 io_oeb[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_75 io_oeb[23] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_42 io_out[28] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_128 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__205__I0 net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_333_ mod.flipflop29.d net1 mod.flipflop29.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_264_ _069_ _072_ _073_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_195_ mod.flipflop8.q _147_ _006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_49_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__290__A1 mod.flipflop36.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_316_ net11 _123_ _124_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_247_ _013_ _016_ _020_ _056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_178_ mod.flipflop33.q _148_ _151_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_6_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__281__A1 _039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_234 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_259 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__250__I _035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__272__A1 mod.flipflop39.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_60 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__263__A1 _134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_281 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__254__A1 _059_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__309__A2 _038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__245__I _050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__155__I _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_207 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_229 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__236__A1 _017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__227__A1 net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__329__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_104 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__160__A3 mod.flipflop36.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_280_ _039_ _060_ _089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_43 io_out[29] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_21 io_out[0] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_54 io_oeb[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_65 io_oeb[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_32 io_out[11] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_17_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_76 io_oeb[24] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__205__I1 net11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_390 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_332_ mod.flipflop29.q net1 mod.flipflop30.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_263_ _134_ _070_ _071_ _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_2
XPHY_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_63 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_74 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_194_ _005_ mod.flipflop12.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_62 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_51 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__290__A2 _058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_315_ _110_ _119_ _122_ _131_ _123_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_246_ _049_ _054_ _055_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_177_ _150_ mod.flipflop37.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__281__A2 _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__272__A2 _080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__362__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__441__I net5 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__263__A2 _070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_229_ mod.flipflop41.q _037_ _038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_2
XFILLER_8_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__254__A2 _062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_219 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__236__A2 _044_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__227__A2 _028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__256__I net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__163__A1 mod.flipflop38.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_116 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__160__A4 mod.flipflop37.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_44 io_out[30] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_55 io_oeb[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_77 io_oeb[25] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_22 io_out[1] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_66 io_oeb[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_33 io_out[12] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_36_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_84 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__205__I2 net12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_391 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_331_ mod.flipflop30.q net1 mod.flipflop31.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_41_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_18_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_64 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_193_ mod.flipflop11.q _147_ _005_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XPHY_86 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_262_ _041_ _052_ _067_ _071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_188 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_75 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__284__B1 _091_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__290__A3 _098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__275__B1 _077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_314_ _142_ _122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_52_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_176_ mod.flipflop36.q _148_ _150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_6_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_245_ _050_ _054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__281__A3 _022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__259__I _134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_239 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_40 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__263__A3 _071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_206 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_261 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_228_ _026_ _036_ _037_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_159_ mod.flipflop40.q _134_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__300__C _108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__311__B _142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__352__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__163__A2 mod.flipflop39.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__182__I _146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_348 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_34 io_out[13] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_23 io_out[2] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_78 io_oeb[26] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_67 io_oeb[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_56 io_oeb[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_45 io_out[31] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_96 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__177__I _150_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__205__I3 net6 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_381 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_370 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_98 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_330_ mod.flipflop32.d net1 mod.flipflop32.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_87 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_43 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_21 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_261_ _055_ _057_ _063_ _070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_41_97 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_192_ _004_ mod.flipflop18.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__293__A1 _054_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__284__A1 mod.flipflop35.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__284__B2 _092_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__275__B2 _056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__275__A1 _061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_85 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_41 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_30 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_244_ _041_ _052_ _053_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_14_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_313_ _121_ mod.flipflop17.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_175_ _149_ mod.flipflop41.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__190__I _003_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_204 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_226 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__257__A1 net4 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__248__A1 _056_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_52 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_227_ net4 _028_ _035_ _036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_273 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_158_ _133_ mod.flipflop8.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__239__B2 _047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__309__B _116_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__311__C _131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__163__A3 mod.flipflop40.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__306__C _047_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__322__B _122_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_24 io_out[3] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_49_416 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_79 io_oeb[27] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_35 io_out[14] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_46 io_out[32] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_57 io_oeb[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_68 io_oeb[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__342__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_393 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_382 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_371 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_99 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_260_ _053_ _064_ _067_ _068_ _069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__365__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__227__B _035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_11 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_33 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_55 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_191_ mod.flipflop14.q _147_ _004_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_41_54 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__293__A2 _062_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__284__A2 _085_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__275__A2 _083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_243_ _049_ _051_ _022_ _052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_53 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_312_ net12 _120_ _121_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_14_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_174_ _134_ _148_ _149_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_6_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_238 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__257__A2 _027_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__193__A1 mod.flipflop11.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__248__A2 _025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_20 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_226_ _030_ _031_ _032_ _034_ _018_ _035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai32_2
X_157_ mod.flipflop33.q _131_ _132_ _133_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_42_285 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__239__A2 net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__166__A1 mod.flipflop19.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__196__I _006_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__157__A1 mod.flipflop33.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_209_ _017_ _018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__320__A1 net10 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__163__A4 mod.flipflop41.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_380 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__311__A1 _110_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_328 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__302__A1 _069_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__322__C _125_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_100 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_25 io_out[4] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_36 io_out[15] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_1_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
Xtiny_user_project_47 io_out[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_58 io_oeb[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_69 io_oeb[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_76 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_177 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_199 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_394 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_383 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_372 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_361 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
X_190_ _003_ mod.flipflop21.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_103 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_67 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_78 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__243__B _022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_280 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_180 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_191 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__332__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__238__B net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_65 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_311_ _110_ _119_ _142_ _131_ _120_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_173_ _147_ _148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_242_ _050_ _051_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__355__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__193__A2 _147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_32 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_225_ _029_ _033_ _034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_8_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_156_ mod.flipflop11.d mod.flipflop8.q _132_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__239__A3 _043_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__166__A2 mod.flipflop20.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__157__A2 _131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_208_ net8 _017_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_24_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_337 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__320__A2 _126_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__311__A2 _119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__302__A2 _072_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xtiny_user_project_26 io_out[5] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_37 io_out[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_48 io_out[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_59 io_oeb[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_39_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_88 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_145 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__296__A1 _058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_167 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_373 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__287__A1 _089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_351 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_35 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_46 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__211__A1 _018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__278__A1 _039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_89 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__269__A1 _028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_292 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_181 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_192 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_22 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_310_ mod.flipflop39.q _111_ _112_ _113_ _118_ _119_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_36_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_172_ _146_ _147_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_241_ _023_ net3 _050_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_218 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__330__D mod.flipflop32.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_44 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_224_ _015_ _033_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_265 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_155_ _130_ _131_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_210 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__325__D mod.flipflop37.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__166__A3 mod.flipflop22.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_207_ _014_ _015_ _016_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__345__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_349 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_139 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__368__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_305 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__262__B _067_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__302__A3 _038_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xtiny_user_project_16 io_oeb[33] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_38 io_out[17] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_27 io_out[6] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_49 io_out[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__296__A2 _098_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_113 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__333__D mod.flipflop29.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_396 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_352 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__287__A2 _083_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_330 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_411 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_25 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__211__A2 _019_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_190 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__278__A2 _075_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__269__A2 _077_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__328__D mod.flipflop34.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_260 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_171 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_182 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_193 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
X_240_ _048_ _049_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_45 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_171_ _135_ _139_ _140_ _145_ _146_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_369_ mod.flipflop38.q net1 mod.flipflop39.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__187__A1 mod.flipflop26.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__178__A1 mod.flipflop33.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_12 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_223_ _018_ _012_ _032_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_42_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__169__A1 mod.flipflop18.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__265__B _028_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_154_ mod.flipflop43.q _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__341__D mod.flipflop21.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__166__A4 mod.flipflop25.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__323__A1 net9 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_206_ net5 net9 net10 net11 mod.flipflop42.q mod.flipflop43.q _015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_30_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__336__D mod.flipflop25.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__305__A1 _070_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__302__A4 _080_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__335__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_17 io_oeb[34] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_39 io_out[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_28 io_out[7] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_29_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_114 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_125 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__358__CLK net15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_397 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_375 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_364 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__202__I _011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_342 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_320 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_331 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_15 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_58 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_47 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_150 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_161 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_183 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_57 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_170_ _141_ _143_ _144_ _145_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_297 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_412 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_368_ mod.flipflop39.q net1 mod.flipflop40.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_299_ _101_ _104_ _108_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__187__A2 _153_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__339__D mod.flipflop22.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_278 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__178__A2 _148_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_24 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_79 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_222_ _019_ _029_ _031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__169__A2 mod.flipflop21.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__281__B _089_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__210__I net7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_315 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_205_ net10 net11 net12 net6 mod.flipflop42.q _130_ _014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_53_329 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__305__A2 _071_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__352__D mod.flipflop5.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_340 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__241__A1 _023_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_189 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__232__A1 _039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__299__A1 _101_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input7_I io_in[18] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_123 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__223__A1 _018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__347__D mod.flipflop12.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
Xtiny_user_project_18 io_oeb[35] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
Xtiny_user_project_29 io_out[8] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_40_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_159 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_310 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_387 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_376 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_365 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_343 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_27 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__325__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__360__D mod.flipflop10.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_162 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_151 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_140 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_173 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_184 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_254 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_240 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_195 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_69 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__279__B _035_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__348__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__234__S _013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_298_ _041_ _082_ _092_ _087_ _062_ _059_ _107_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_367_ mod.flipflop41.d net1 mod.flipflop41.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_9_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__355__D mod.flipflop2.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_36 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_257 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_224 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__169__A3 mod.flipflop23.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_221_ _019_ _029_ _030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_18_243 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_202 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_327 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__276__C _084_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_204_ _012_ _013_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__241__A2 net3 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__287__B _065_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_341 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__232__A2 _040_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__299__A2 _104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_157 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__223__A2 _012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__363__D mod.flipflop1.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
Xtiny_user_project_19 io_oeb[36] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_44_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_366 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_355 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_300 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_322 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_403 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_399 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__358__D mod.flipflop16.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_119 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_160 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_7 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__284__C mod.flipflop34.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__199__A1 _007_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_8 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_270 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_252 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_230 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_163 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_174 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_185 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_196 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_299 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_277 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_244 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_37 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_26 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_318 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_414 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_366_ mod.flipflop41.q net1 mod.flipflop42.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_13_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_297_ _101_ _104_ _105_ _106_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__314__I _142_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_81 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_211 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_222 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_258 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__224__I _015_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_220_ _014_ _029_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_269 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__169__A4 mod.flipflop24.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_80 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_349_ mod.flipflop9.d net1 mod.flipflop11.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__366__D mod.flipflop41.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__308__A1 _026_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__338__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_339 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
X_203_ net9 net10 net11 net12 mod.flipflop42.q _130_ _012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_7_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_317 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__226__B1 _034_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_309 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_353 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_283 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_350 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_147 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__289__I0 _095_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_117 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_378 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_367 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_345 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_334 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_301 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_312 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_323 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_39 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_194 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_209 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__199__A2 _008_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_282 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_242 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_172 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__369__D mod.flipflop38.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_264 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_164 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_153 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_142 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_131 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_120 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_175 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_186 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_197 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_49 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__295__C _058_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_245 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_296_ _058_ _098_ mod.flipflop36.q _105_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_365_ mod.flipflop42.q net1 mod.flipflop43.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_45_289 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__280__A1 _039_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__271__A1 _022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_16 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_237 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_101 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__262__A1 _041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_93 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_92 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_70 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_279_ _040_ _061_ _035_ _088_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_348_ mod.flipflop11.d net1 mod.flipflop11.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_392 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__253__A1 _060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__308__A2 _036_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_307 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__244__A1 _041_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_215 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_202_ _011_ mod.flipflop2.d vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_output14_I net14 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__235__A1 _012_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_384 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_332 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__226__A1 _030_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__226__B2 _018_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__217__A1 _022_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_115 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__328__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_409 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_354 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_170 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__289__I1 _097_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_129 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_368 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_346 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_335 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_413 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input5_I io_in[16] vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_302 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_19 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_45_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__203__S0 mod.flipflop42.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_132 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_110 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_121 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_165 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_154 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_143 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_187 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_198 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_405 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_17 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_176 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
X_295_ _082_ _102_ _103_ _058_ _104_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_364_ mod.flipflop1.d net1 mod.flipflop1.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_61 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__280__A2 _060_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_66 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_408 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_246 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_28 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__271__A2 _074_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_419 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_279 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_293 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_179 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_389 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__262__A2 _052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__361__CLK net1 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_347_ mod.flipflop12.d net1 mod.flipflop12.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_278_ _039_ _075_ _087_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_271 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_360 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__253__A2 _061_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__251__I net2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_319 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__244__A2 _052_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
X_201_ net15 _010_ _011_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__180__A1 mod.flipflop32.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__235__A2 _014_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_208 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__171__A1 _135_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_344 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__226__A2 _031_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_18 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_388 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__162__A1 mod.flipflop26.q vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__217__A2 _025_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_385 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_212 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_105 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_127 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_31 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_50 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_73 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_303 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_369 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_347 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_2 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_108 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_325 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_314 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_130 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_152 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_417 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_141 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__203__S1 _130_ vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_166 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_155 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_144 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_133 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_111 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_122 vccd1 vssd1 gf180mcu_fd_sc_mcu7t5v0__filltie
.ends

