magic
tech gf180mcuC
magscale 1 10
timestamp 1669308287
<< metal1 >>
rect 25554 48974 25566 49026
rect 25618 49023 25630 49026
rect 26450 49023 26462 49026
rect 25618 48977 26462 49023
rect 25618 48974 25630 48977
rect 26450 48974 26462 48977
rect 26514 48974 26526 49026
rect 22978 48750 22990 48802
rect 23042 48799 23054 48802
rect 27010 48799 27022 48802
rect 23042 48753 27022 48799
rect 23042 48750 23054 48753
rect 27010 48750 27022 48753
rect 27074 48750 27086 48802
rect 23650 47742 23662 47794
rect 23714 47791 23726 47794
rect 23986 47791 23998 47794
rect 23714 47745 23998 47791
rect 23714 47742 23726 47745
rect 23986 47742 23998 47745
rect 24050 47791 24062 47794
rect 27010 47791 27022 47794
rect 24050 47745 27022 47791
rect 24050 47742 24062 47745
rect 27010 47742 27022 47745
rect 27074 47742 27086 47794
rect 13906 47406 13918 47458
rect 13970 47455 13982 47458
rect 15474 47455 15486 47458
rect 13970 47409 15486 47455
rect 13970 47406 13982 47409
rect 15474 47406 15486 47409
rect 15538 47455 15550 47458
rect 16706 47455 16718 47458
rect 15538 47409 16718 47455
rect 15538 47406 15550 47409
rect 16706 47406 16718 47409
rect 16770 47406 16782 47458
rect 14690 47182 14702 47234
rect 14754 47231 14766 47234
rect 16034 47231 16046 47234
rect 14754 47185 16046 47231
rect 14754 47182 14766 47185
rect 16034 47182 16046 47185
rect 16098 47182 16110 47234
rect 8306 46958 8318 47010
rect 8370 47007 8382 47010
rect 8530 47007 8542 47010
rect 8370 46961 8542 47007
rect 8370 46958 8382 46961
rect 8530 46958 8542 46961
rect 8594 46958 8606 47010
rect 32274 46734 32286 46786
rect 32338 46783 32350 46786
rect 33394 46783 33406 46786
rect 32338 46737 33406 46783
rect 32338 46734 32350 46737
rect 33394 46734 33406 46737
rect 33458 46734 33470 46786
rect 27682 46510 27694 46562
rect 27746 46559 27758 46562
rect 29810 46559 29822 46562
rect 27746 46513 29822 46559
rect 27746 46510 27758 46513
rect 29810 46510 29822 46513
rect 29874 46559 29886 46562
rect 31938 46559 31950 46562
rect 29874 46513 31950 46559
rect 29874 46510 29886 46513
rect 31938 46510 31950 46513
rect 32002 46510 32014 46562
rect 2034 46398 2046 46450
rect 2098 46447 2110 46450
rect 2706 46447 2718 46450
rect 2098 46401 2718 46447
rect 2098 46398 2110 46401
rect 2706 46398 2718 46401
rect 2770 46398 2782 46450
rect 8866 46398 8878 46450
rect 8930 46447 8942 46450
rect 9426 46447 9438 46450
rect 8930 46401 9438 46447
rect 8930 46398 8942 46401
rect 9426 46398 9438 46401
rect 9490 46398 9502 46450
rect 1344 46282 48608 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 48608 46282
rect 1344 46196 48608 46230
rect 28366 46114 28418 46126
rect 28366 46050 28418 46062
rect 5854 46002 5906 46014
rect 4050 45950 4062 46002
rect 4114 45950 4126 46002
rect 5854 45938 5906 45950
rect 7198 46002 7250 46014
rect 7198 45938 7250 45950
rect 9774 46002 9826 46014
rect 26350 46002 26402 46014
rect 38446 46002 38498 46014
rect 11890 45950 11902 46002
rect 11954 45950 11966 46002
rect 17714 45950 17726 46002
rect 17778 45950 17790 46002
rect 19842 45950 19854 46002
rect 19906 45950 19918 46002
rect 22194 45950 22206 46002
rect 22258 45950 22270 46002
rect 24322 45950 24334 46002
rect 24386 45950 24398 46002
rect 25778 45950 25790 46002
rect 25842 45950 25854 46002
rect 33394 45950 33406 46002
rect 33458 45950 33470 46002
rect 35634 45950 35646 46002
rect 35698 45950 35710 46002
rect 9774 45938 9826 45950
rect 26350 45938 26402 45950
rect 38446 45938 38498 45950
rect 38894 46002 38946 46014
rect 38894 45938 38946 45950
rect 39342 46002 39394 46014
rect 39342 45938 39394 45950
rect 1822 45890 1874 45902
rect 27806 45890 27858 45902
rect 41806 45890 41858 45902
rect 4834 45838 4846 45890
rect 4898 45838 4910 45890
rect 13570 45838 13582 45890
rect 13634 45838 13646 45890
rect 20626 45838 20638 45890
rect 20690 45838 20702 45890
rect 21522 45838 21534 45890
rect 21586 45838 21598 45890
rect 26002 45838 26014 45890
rect 26066 45838 26078 45890
rect 34178 45838 34190 45890
rect 34242 45838 34254 45890
rect 36082 45838 36094 45890
rect 36146 45838 36158 45890
rect 1822 45826 1874 45838
rect 27806 45826 27858 45838
rect 41806 45826 41858 45838
rect 2158 45778 2210 45790
rect 2158 45714 2210 45726
rect 2718 45778 2770 45790
rect 2718 45714 2770 45726
rect 7646 45778 7698 45790
rect 7646 45714 7698 45726
rect 8878 45778 8930 45790
rect 8878 45714 8930 45726
rect 10334 45778 10386 45790
rect 10334 45714 10386 45726
rect 11006 45778 11058 45790
rect 11006 45714 11058 45726
rect 11566 45778 11618 45790
rect 11566 45714 11618 45726
rect 12462 45778 12514 45790
rect 27470 45778 27522 45790
rect 15362 45726 15374 45778
rect 15426 45726 15438 45778
rect 27346 45726 27358 45778
rect 27410 45726 27422 45778
rect 12462 45714 12514 45726
rect 27470 45714 27522 45726
rect 27582 45778 27634 45790
rect 27582 45714 27634 45726
rect 28478 45778 28530 45790
rect 28478 45714 28530 45726
rect 30158 45778 30210 45790
rect 30158 45714 30210 45726
rect 31502 45778 31554 45790
rect 31502 45714 31554 45726
rect 32062 45778 32114 45790
rect 32062 45714 32114 45726
rect 37886 45778 37938 45790
rect 37886 45714 37938 45726
rect 39902 45778 39954 45790
rect 39902 45714 39954 45726
rect 41358 45778 41410 45790
rect 41358 45714 41410 45726
rect 43262 45778 43314 45790
rect 43262 45714 43314 45726
rect 48078 45778 48130 45790
rect 48078 45714 48130 45726
rect 6190 45666 6242 45678
rect 6190 45602 6242 45614
rect 6638 45666 6690 45678
rect 6638 45602 6690 45614
rect 8206 45666 8258 45678
rect 8206 45602 8258 45614
rect 11790 45666 11842 45678
rect 11790 45602 11842 45614
rect 12798 45666 12850 45678
rect 12798 45602 12850 45614
rect 16718 45666 16770 45678
rect 16718 45602 16770 45614
rect 27694 45666 27746 45678
rect 29598 45666 29650 45678
rect 29250 45614 29262 45666
rect 29314 45614 29326 45666
rect 27694 45602 27746 45614
rect 29598 45602 29650 45614
rect 31166 45666 31218 45678
rect 31166 45602 31218 45614
rect 37102 45666 37154 45678
rect 37102 45602 37154 45614
rect 40910 45666 40962 45678
rect 40910 45602 40962 45614
rect 1344 45498 48608 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 48608 45498
rect 1344 45412 48608 45446
rect 1822 45330 1874 45342
rect 1822 45266 1874 45278
rect 2494 45330 2546 45342
rect 2494 45266 2546 45278
rect 3166 45330 3218 45342
rect 3166 45266 3218 45278
rect 4622 45330 4674 45342
rect 4622 45266 4674 45278
rect 5070 45330 5122 45342
rect 5070 45266 5122 45278
rect 5966 45330 6018 45342
rect 5966 45266 6018 45278
rect 8206 45330 8258 45342
rect 8206 45266 8258 45278
rect 8542 45330 8594 45342
rect 8542 45266 8594 45278
rect 9102 45330 9154 45342
rect 9102 45266 9154 45278
rect 10670 45330 10722 45342
rect 10670 45266 10722 45278
rect 12238 45330 12290 45342
rect 12238 45266 12290 45278
rect 31502 45330 31554 45342
rect 31502 45266 31554 45278
rect 32062 45330 32114 45342
rect 32062 45266 32114 45278
rect 32398 45330 32450 45342
rect 32398 45266 32450 45278
rect 36206 45330 36258 45342
rect 36206 45266 36258 45278
rect 37102 45330 37154 45342
rect 37102 45266 37154 45278
rect 38446 45330 38498 45342
rect 38446 45266 38498 45278
rect 39342 45330 39394 45342
rect 39342 45266 39394 45278
rect 39790 45330 39842 45342
rect 39790 45266 39842 45278
rect 40686 45330 40738 45342
rect 40686 45266 40738 45278
rect 11118 45218 11170 45230
rect 11118 45154 11170 45166
rect 11454 45218 11506 45230
rect 11454 45154 11506 45166
rect 13470 45218 13522 45230
rect 28030 45218 28082 45230
rect 18610 45166 18622 45218
rect 18674 45166 18686 45218
rect 22978 45166 22990 45218
rect 23042 45166 23054 45218
rect 26002 45166 26014 45218
rect 26066 45166 26078 45218
rect 13470 45154 13522 45166
rect 28030 45154 28082 45166
rect 28926 45218 28978 45230
rect 28926 45154 28978 45166
rect 29262 45218 29314 45230
rect 29262 45154 29314 45166
rect 30382 45218 30434 45230
rect 30382 45154 30434 45166
rect 34862 45218 34914 45230
rect 34862 45154 34914 45166
rect 6750 45106 6802 45118
rect 6750 45042 6802 45054
rect 13246 45106 13298 45118
rect 24446 45106 24498 45118
rect 26574 45106 26626 45118
rect 14018 45054 14030 45106
rect 14082 45054 14094 45106
rect 17714 45054 17726 45106
rect 17778 45054 17790 45106
rect 19506 45054 19518 45106
rect 19570 45054 19582 45106
rect 23090 45054 23102 45106
rect 23154 45054 23166 45106
rect 23762 45054 23774 45106
rect 23826 45054 23838 45106
rect 25778 45054 25790 45106
rect 25842 45054 25854 45106
rect 13246 45042 13298 45054
rect 24446 45042 24498 45054
rect 26574 45042 26626 45054
rect 28142 45106 28194 45118
rect 29374 45106 29426 45118
rect 33630 45106 33682 45118
rect 28354 45054 28366 45106
rect 28418 45054 28430 45106
rect 30034 45054 30046 45106
rect 30098 45054 30110 45106
rect 28142 45042 28194 45054
rect 29374 45042 29426 45054
rect 33630 45042 33682 45054
rect 4174 44994 4226 45006
rect 4174 44930 4226 44942
rect 5518 44994 5570 45006
rect 5518 44930 5570 44942
rect 6302 44994 6354 45006
rect 6302 44930 6354 44942
rect 7310 44994 7362 45006
rect 7310 44930 7362 44942
rect 7758 44994 7810 45006
rect 7758 44930 7810 44942
rect 9774 44994 9826 45006
rect 9774 44930 9826 44942
rect 10222 44994 10274 45006
rect 10222 44930 10274 44942
rect 12910 44994 12962 45006
rect 24894 44994 24946 45006
rect 29038 44994 29090 45006
rect 14802 44942 14814 44994
rect 14866 44942 14878 44994
rect 16930 44942 16942 44994
rect 16994 44942 17006 44994
rect 20290 44942 20302 44994
rect 20354 44942 20366 44994
rect 22418 44942 22430 44994
rect 22482 44942 22494 44994
rect 27570 44942 27582 44994
rect 27634 44942 27646 44994
rect 12910 44930 12962 44942
rect 24894 44930 24946 44942
rect 29038 44930 29090 44942
rect 31054 44994 31106 45006
rect 31054 44930 31106 44942
rect 32846 44994 32898 45006
rect 32846 44930 32898 44942
rect 33966 44994 34018 45006
rect 33966 44930 34018 44942
rect 34414 44994 34466 45006
rect 34414 44930 34466 44942
rect 35310 44994 35362 45006
rect 35310 44930 35362 44942
rect 35758 44994 35810 45006
rect 35758 44930 35810 44942
rect 36654 44994 36706 45006
rect 36654 44930 36706 44942
rect 37550 44994 37602 45006
rect 37550 44930 37602 44942
rect 37998 44994 38050 45006
rect 37998 44930 38050 44942
rect 38894 44994 38946 45006
rect 38894 44930 38946 44942
rect 40238 44994 40290 45006
rect 40238 44930 40290 44942
rect 12014 44882 12066 44894
rect 12014 44818 12066 44830
rect 12350 44882 12402 44894
rect 12350 44818 12402 44830
rect 24558 44882 24610 44894
rect 24558 44818 24610 44830
rect 26910 44882 26962 44894
rect 26910 44818 26962 44830
rect 30046 44882 30098 44894
rect 30046 44818 30098 44830
rect 30942 44882 30994 44894
rect 31938 44830 31950 44882
rect 32002 44879 32014 44882
rect 32834 44879 32846 44882
rect 32002 44833 32846 44879
rect 32002 44830 32014 44833
rect 32834 44830 32846 44833
rect 32898 44830 32910 44882
rect 36978 44830 36990 44882
rect 37042 44879 37054 44882
rect 37986 44879 37998 44882
rect 37042 44833 37998 44879
rect 37042 44830 37054 44833
rect 37986 44830 37998 44833
rect 38050 44830 38062 44882
rect 30942 44818 30994 44830
rect 1344 44714 48608 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 48608 44714
rect 1344 44628 48608 44662
rect 11454 44546 11506 44558
rect 11454 44482 11506 44494
rect 11790 44546 11842 44558
rect 11790 44482 11842 44494
rect 28702 44546 28754 44558
rect 33954 44494 33966 44546
rect 34018 44543 34030 44546
rect 34626 44543 34638 44546
rect 34018 44497 34638 44543
rect 34018 44494 34030 44497
rect 34626 44494 34638 44497
rect 34690 44494 34702 44546
rect 28702 44482 28754 44494
rect 3726 44434 3778 44446
rect 3726 44370 3778 44382
rect 4174 44434 4226 44446
rect 4174 44370 4226 44382
rect 5070 44434 5122 44446
rect 5070 44370 5122 44382
rect 6750 44434 6802 44446
rect 6750 44370 6802 44382
rect 7198 44434 7250 44446
rect 7198 44370 7250 44382
rect 8094 44434 8146 44446
rect 8094 44370 8146 44382
rect 9774 44434 9826 44446
rect 9774 44370 9826 44382
rect 11230 44434 11282 44446
rect 31166 44434 31218 44446
rect 15250 44382 15262 44434
rect 15314 44382 15326 44434
rect 17378 44382 17390 44434
rect 17442 44382 17454 44434
rect 18722 44382 18734 44434
rect 18786 44382 18798 44434
rect 20850 44382 20862 44434
rect 20914 44382 20926 44434
rect 22418 44382 22430 44434
rect 22482 44382 22494 44434
rect 24546 44382 24558 44434
rect 24610 44382 24622 44434
rect 25890 44382 25902 44434
rect 25954 44382 25966 44434
rect 28018 44382 28030 44434
rect 28082 44382 28094 44434
rect 11230 44370 11282 44382
rect 31166 44370 31218 44382
rect 33070 44434 33122 44446
rect 33070 44370 33122 44382
rect 33966 44434 34018 44446
rect 33966 44370 34018 44382
rect 37438 44434 37490 44446
rect 37438 44370 37490 44382
rect 38334 44434 38386 44446
rect 38334 44370 38386 44382
rect 39678 44434 39730 44446
rect 39678 44370 39730 44382
rect 4622 44322 4674 44334
rect 12350 44322 12402 44334
rect 3042 44270 3054 44322
rect 3106 44270 3118 44322
rect 10434 44270 10446 44322
rect 10498 44270 10510 44322
rect 4622 44258 4674 44270
rect 12350 44258 12402 44270
rect 12910 44322 12962 44334
rect 12910 44258 12962 44270
rect 14030 44322 14082 44334
rect 29822 44322 29874 44334
rect 31054 44322 31106 44334
rect 14466 44270 14478 44322
rect 14530 44270 14542 44322
rect 17938 44270 17950 44322
rect 18002 44270 18014 44322
rect 21634 44270 21646 44322
rect 21698 44270 21710 44322
rect 25218 44270 25230 44322
rect 25282 44270 25294 44322
rect 30706 44270 30718 44322
rect 30770 44270 30782 44322
rect 14030 44258 14082 44270
rect 29822 44258 29874 44270
rect 31054 44258 31106 44270
rect 31838 44322 31890 44334
rect 31838 44258 31890 44270
rect 38782 44322 38834 44334
rect 38782 44258 38834 44270
rect 5854 44210 5906 44222
rect 2146 44158 2158 44210
rect 2210 44158 2222 44210
rect 5854 44146 5906 44158
rect 10670 44210 10722 44222
rect 10670 44146 10722 44158
rect 12574 44210 12626 44222
rect 12574 44146 12626 44158
rect 13694 44210 13746 44222
rect 13694 44146 13746 44158
rect 13806 44210 13858 44222
rect 13806 44146 13858 44158
rect 28702 44210 28754 44222
rect 28702 44146 28754 44158
rect 28814 44210 28866 44222
rect 35310 44210 35362 44222
rect 32162 44158 32174 44210
rect 32226 44158 32238 44210
rect 28814 44146 28866 44158
rect 35310 44146 35362 44158
rect 6190 44098 6242 44110
rect 6190 44034 6242 44046
rect 7646 44098 7698 44110
rect 7646 44034 7698 44046
rect 8430 44098 8482 44110
rect 8430 44034 8482 44046
rect 8990 44098 9042 44110
rect 8990 44034 9042 44046
rect 9438 44098 9490 44110
rect 9438 44034 9490 44046
rect 12686 44098 12738 44110
rect 12686 44034 12738 44046
rect 29598 44098 29650 44110
rect 29598 44034 29650 44046
rect 29710 44098 29762 44110
rect 29710 44034 29762 44046
rect 30046 44098 30098 44110
rect 30046 44034 30098 44046
rect 31278 44098 31330 44110
rect 31278 44034 31330 44046
rect 32734 44098 32786 44110
rect 32734 44034 32786 44046
rect 33518 44098 33570 44110
rect 33518 44034 33570 44046
rect 34526 44098 34578 44110
rect 34526 44034 34578 44046
rect 34974 44098 35026 44110
rect 34974 44034 35026 44046
rect 35758 44098 35810 44110
rect 35758 44034 35810 44046
rect 36206 44098 36258 44110
rect 36206 44034 36258 44046
rect 36654 44098 36706 44110
rect 36654 44034 36706 44046
rect 37886 44098 37938 44110
rect 37886 44034 37938 44046
rect 39230 44098 39282 44110
rect 39230 44034 39282 44046
rect 40126 44098 40178 44110
rect 40126 44034 40178 44046
rect 1344 43930 48608 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 48608 43930
rect 1344 43844 48608 43878
rect 1934 43762 1986 43774
rect 1934 43698 1986 43710
rect 10670 43762 10722 43774
rect 10670 43698 10722 43710
rect 11678 43762 11730 43774
rect 11678 43698 11730 43710
rect 18958 43762 19010 43774
rect 18958 43698 19010 43710
rect 31054 43762 31106 43774
rect 31054 43698 31106 43710
rect 31726 43762 31778 43774
rect 31726 43698 31778 43710
rect 37102 43762 37154 43774
rect 37102 43698 37154 43710
rect 38894 43762 38946 43774
rect 38894 43698 38946 43710
rect 40686 43762 40738 43774
rect 40686 43698 40738 43710
rect 47742 43762 47794 43774
rect 47742 43698 47794 43710
rect 3726 43650 3778 43662
rect 3726 43586 3778 43598
rect 4958 43650 5010 43662
rect 4958 43586 5010 43598
rect 8206 43650 8258 43662
rect 8206 43586 8258 43598
rect 9886 43650 9938 43662
rect 9886 43586 9938 43598
rect 11454 43650 11506 43662
rect 11454 43586 11506 43598
rect 11790 43650 11842 43662
rect 31838 43650 31890 43662
rect 14802 43598 14814 43650
rect 14866 43598 14878 43650
rect 17938 43598 17950 43650
rect 18002 43598 18014 43650
rect 18386 43598 18398 43650
rect 18450 43598 18462 43650
rect 27794 43598 27806 43650
rect 27858 43598 27870 43650
rect 11790 43586 11842 43598
rect 31838 43586 31890 43598
rect 32062 43650 32114 43662
rect 32062 43586 32114 43598
rect 33966 43650 34018 43662
rect 33966 43586 34018 43598
rect 4174 43538 4226 43550
rect 4174 43474 4226 43486
rect 6750 43538 6802 43550
rect 11230 43538 11282 43550
rect 13470 43538 13522 43550
rect 18622 43538 18674 43550
rect 24110 43538 24162 43550
rect 29710 43538 29762 43550
rect 10434 43486 10446 43538
rect 10498 43486 10510 43538
rect 13010 43486 13022 43538
rect 13074 43486 13086 43538
rect 14018 43486 14030 43538
rect 14082 43486 14094 43538
rect 19618 43486 19630 43538
rect 19682 43486 19694 43538
rect 23314 43486 23326 43538
rect 23378 43486 23390 43538
rect 24546 43486 24558 43538
rect 24610 43486 24622 43538
rect 28466 43486 28478 43538
rect 28530 43486 28542 43538
rect 29474 43486 29486 43538
rect 29538 43486 29550 43538
rect 6750 43474 6802 43486
rect 11230 43474 11282 43486
rect 13470 43474 13522 43486
rect 18622 43474 18674 43486
rect 24110 43474 24162 43486
rect 29710 43474 29762 43486
rect 29822 43538 29874 43550
rect 29822 43474 29874 43486
rect 30046 43538 30098 43550
rect 30046 43474 30098 43486
rect 30718 43538 30770 43550
rect 30718 43474 30770 43486
rect 30830 43538 30882 43550
rect 30830 43474 30882 43486
rect 30942 43538 30994 43550
rect 32398 43538 32450 43550
rect 31266 43486 31278 43538
rect 31330 43486 31342 43538
rect 30942 43474 30994 43486
rect 32398 43474 32450 43486
rect 37998 43538 38050 43550
rect 37998 43474 38050 43486
rect 48078 43538 48130 43550
rect 48078 43474 48130 43486
rect 2382 43426 2434 43438
rect 2382 43362 2434 43374
rect 2830 43426 2882 43438
rect 2830 43362 2882 43374
rect 3166 43426 3218 43438
rect 3166 43362 3218 43374
rect 4622 43426 4674 43438
rect 4622 43362 4674 43374
rect 5518 43426 5570 43438
rect 5518 43362 5570 43374
rect 5966 43426 6018 43438
rect 5966 43362 6018 43374
rect 6302 43426 6354 43438
rect 6302 43362 6354 43374
rect 7310 43426 7362 43438
rect 7310 43362 7362 43374
rect 7758 43426 7810 43438
rect 7758 43362 7810 43374
rect 8654 43426 8706 43438
rect 8654 43362 8706 43374
rect 9102 43426 9154 43438
rect 29038 43426 29090 43438
rect 12674 43374 12686 43426
rect 12738 43374 12750 43426
rect 16930 43374 16942 43426
rect 16994 43374 17006 43426
rect 20402 43374 20414 43426
rect 20466 43374 20478 43426
rect 22530 43374 22542 43426
rect 22594 43374 22606 43426
rect 23650 43374 23662 43426
rect 23714 43374 23726 43426
rect 25666 43374 25678 43426
rect 25730 43374 25742 43426
rect 9102 43362 9154 43374
rect 29038 43362 29090 43374
rect 32734 43426 32786 43438
rect 32734 43362 32786 43374
rect 33518 43426 33570 43438
rect 33518 43362 33570 43374
rect 34414 43426 34466 43438
rect 34414 43362 34466 43374
rect 34862 43426 34914 43438
rect 34862 43362 34914 43374
rect 35310 43426 35362 43438
rect 35310 43362 35362 43374
rect 35758 43426 35810 43438
rect 35758 43362 35810 43374
rect 36206 43426 36258 43438
rect 36206 43362 36258 43374
rect 36654 43426 36706 43438
rect 36654 43362 36706 43374
rect 37550 43426 37602 43438
rect 37550 43362 37602 43374
rect 38446 43426 38498 43438
rect 38446 43362 38498 43374
rect 39342 43426 39394 43438
rect 39342 43362 39394 43374
rect 39790 43426 39842 43438
rect 39790 43362 39842 43374
rect 40238 43426 40290 43438
rect 40238 43362 40290 43374
rect 47294 43426 47346 43438
rect 47294 43362 47346 43374
rect 6962 43262 6974 43314
rect 7026 43311 7038 43314
rect 7746 43311 7758 43314
rect 7026 43265 7758 43311
rect 7026 43262 7038 43265
rect 7746 43262 7758 43265
rect 7810 43262 7822 43314
rect 23538 43262 23550 43314
rect 23602 43262 23614 43314
rect 34178 43262 34190 43314
rect 34242 43311 34254 43314
rect 35410 43311 35422 43314
rect 34242 43265 35422 43311
rect 34242 43262 34254 43265
rect 35410 43262 35422 43265
rect 35474 43262 35486 43314
rect 1344 43146 48608 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 48608 43146
rect 1344 43060 48608 43094
rect 28702 42978 28754 42990
rect 28702 42914 28754 42926
rect 29934 42978 29986 42990
rect 29934 42914 29986 42926
rect 30382 42978 30434 42990
rect 34514 42926 34526 42978
rect 34578 42975 34590 42978
rect 34578 42929 35583 42975
rect 34578 42926 34590 42929
rect 30382 42914 30434 42926
rect 2830 42866 2882 42878
rect 2830 42802 2882 42814
rect 3278 42866 3330 42878
rect 3278 42802 3330 42814
rect 7310 42866 7362 42878
rect 30158 42866 30210 42878
rect 9986 42814 9998 42866
rect 10050 42814 10062 42866
rect 15250 42814 15262 42866
rect 15314 42814 15326 42866
rect 17378 42814 17390 42866
rect 17442 42814 17454 42866
rect 20850 42814 20862 42866
rect 20914 42814 20926 42866
rect 21634 42814 21646 42866
rect 21698 42814 21710 42866
rect 23762 42814 23774 42866
rect 23826 42814 23838 42866
rect 25106 42814 25118 42866
rect 25170 42814 25182 42866
rect 27234 42814 27246 42866
rect 27298 42814 27310 42866
rect 7310 42802 7362 42814
rect 30158 42802 30210 42814
rect 30606 42866 30658 42878
rect 30606 42802 30658 42814
rect 34414 42866 34466 42878
rect 34414 42802 34466 42814
rect 4174 42754 4226 42766
rect 13694 42754 13746 42766
rect 12898 42702 12910 42754
rect 12962 42702 12974 42754
rect 4174 42690 4226 42702
rect 13694 42690 13746 42702
rect 14030 42754 14082 42766
rect 28590 42754 28642 42766
rect 14466 42702 14478 42754
rect 14530 42702 14542 42754
rect 17938 42702 17950 42754
rect 18002 42702 18014 42754
rect 24546 42702 24558 42754
rect 24610 42702 24622 42754
rect 27906 42702 27918 42754
rect 27970 42702 27982 42754
rect 14030 42690 14082 42702
rect 28590 42690 28642 42702
rect 32846 42754 32898 42766
rect 32846 42690 32898 42702
rect 8206 42642 8258 42654
rect 8206 42578 8258 42590
rect 9102 42642 9154 42654
rect 31390 42642 31442 42654
rect 12114 42590 12126 42642
rect 12178 42590 12190 42642
rect 18722 42590 18734 42642
rect 18786 42590 18798 42642
rect 9102 42578 9154 42590
rect 31390 42578 31442 42590
rect 31502 42642 31554 42654
rect 33070 42642 33122 42654
rect 31602 42590 31614 42642
rect 31666 42590 31678 42642
rect 31502 42578 31554 42590
rect 33070 42578 33122 42590
rect 33742 42642 33794 42654
rect 33742 42578 33794 42590
rect 33966 42642 34018 42654
rect 33966 42578 34018 42590
rect 1822 42530 1874 42542
rect 1822 42466 1874 42478
rect 3726 42530 3778 42542
rect 3726 42466 3778 42478
rect 4622 42530 4674 42542
rect 4622 42466 4674 42478
rect 5070 42530 5122 42542
rect 5070 42466 5122 42478
rect 5854 42530 5906 42542
rect 5854 42466 5906 42478
rect 6302 42530 6354 42542
rect 6302 42466 6354 42478
rect 6750 42530 6802 42542
rect 6750 42466 6802 42478
rect 7758 42530 7810 42542
rect 7758 42466 7810 42478
rect 8542 42530 8594 42542
rect 8542 42466 8594 42478
rect 9214 42530 9266 42542
rect 9214 42466 9266 42478
rect 9326 42530 9378 42542
rect 9326 42466 9378 42478
rect 13806 42530 13858 42542
rect 13806 42466 13858 42478
rect 28702 42530 28754 42542
rect 28702 42466 28754 42478
rect 29486 42530 29538 42542
rect 29486 42466 29538 42478
rect 31166 42530 31218 42542
rect 31166 42466 31218 42478
rect 31278 42530 31330 42542
rect 33854 42530 33906 42542
rect 32498 42478 32510 42530
rect 32562 42478 32574 42530
rect 31278 42466 31330 42478
rect 33854 42466 33906 42478
rect 34862 42530 34914 42542
rect 34862 42466 34914 42478
rect 35310 42530 35362 42542
rect 35537 42527 35583 42929
rect 36206 42866 36258 42878
rect 36206 42802 36258 42814
rect 37998 42866 38050 42878
rect 37998 42802 38050 42814
rect 35758 42754 35810 42766
rect 35758 42690 35810 42702
rect 36654 42754 36706 42766
rect 36654 42690 36706 42702
rect 40126 42642 40178 42654
rect 40126 42578 40178 42590
rect 37438 42530 37490 42542
rect 35634 42527 35646 42530
rect 35537 42481 35646 42527
rect 35634 42478 35646 42481
rect 35698 42478 35710 42530
rect 35310 42466 35362 42478
rect 37438 42466 37490 42478
rect 38446 42530 38498 42542
rect 38446 42466 38498 42478
rect 38782 42530 38834 42542
rect 38782 42466 38834 42478
rect 39230 42530 39282 42542
rect 39230 42466 39282 42478
rect 39678 42530 39730 42542
rect 39678 42466 39730 42478
rect 40574 42530 40626 42542
rect 40574 42466 40626 42478
rect 1344 42362 48608 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 48608 42362
rect 1344 42276 48608 42310
rect 18286 42194 18338 42206
rect 18286 42130 18338 42142
rect 34974 42194 35026 42206
rect 34974 42130 35026 42142
rect 36878 42194 36930 42206
rect 36878 42130 36930 42142
rect 38222 42194 38274 42206
rect 38222 42130 38274 42142
rect 6974 42082 7026 42094
rect 6974 42018 7026 42030
rect 7534 42082 7586 42094
rect 7534 42018 7586 42030
rect 7870 42082 7922 42094
rect 7870 42018 7922 42030
rect 8430 42082 8482 42094
rect 8430 42018 8482 42030
rect 8990 42082 9042 42094
rect 8990 42018 9042 42030
rect 9886 42082 9938 42094
rect 9886 42018 9938 42030
rect 9998 42082 10050 42094
rect 9998 42018 10050 42030
rect 22766 42082 22818 42094
rect 22766 42018 22818 42030
rect 31950 42082 32002 42094
rect 31950 42018 32002 42030
rect 34862 42082 34914 42094
rect 34862 42018 34914 42030
rect 2158 41970 2210 41982
rect 2158 41906 2210 41918
rect 5182 41970 5234 41982
rect 5182 41906 5234 41918
rect 5742 41970 5794 41982
rect 5742 41906 5794 41918
rect 6638 41970 6690 41982
rect 6638 41906 6690 41918
rect 8654 41970 8706 41982
rect 17838 41970 17890 41982
rect 10546 41918 10558 41970
rect 10610 41918 10622 41970
rect 14130 41918 14142 41970
rect 14194 41918 14206 41970
rect 14802 41918 14814 41970
rect 14866 41918 14878 41970
rect 8654 41906 8706 41918
rect 17838 41906 17890 41918
rect 18398 41970 18450 41982
rect 24110 41970 24162 41982
rect 22082 41918 22094 41970
rect 22146 41918 22158 41970
rect 18398 41906 18450 41918
rect 24110 41906 24162 41918
rect 24334 41970 24386 41982
rect 30046 41970 30098 41982
rect 34190 41970 34242 41982
rect 25778 41918 25790 41970
rect 25842 41918 25854 41970
rect 29810 41918 29822 41970
rect 29874 41918 29886 41970
rect 30370 41918 30382 41970
rect 30434 41918 30446 41970
rect 30706 41918 30718 41970
rect 30770 41918 30782 41970
rect 24334 41906 24386 41918
rect 30046 41906 30098 41918
rect 34190 41906 34242 41918
rect 37326 41970 37378 41982
rect 37326 41906 37378 41918
rect 37774 41970 37826 41982
rect 37774 41906 37826 41918
rect 2606 41858 2658 41870
rect 2606 41794 2658 41806
rect 3054 41858 3106 41870
rect 3054 41794 3106 41806
rect 3502 41858 3554 41870
rect 3502 41794 3554 41806
rect 3950 41858 4002 41870
rect 3950 41794 4002 41806
rect 4398 41858 4450 41870
rect 4398 41794 4450 41806
rect 4846 41858 4898 41870
rect 4846 41794 4898 41806
rect 6078 41858 6130 41870
rect 6078 41794 6130 41806
rect 8878 41858 8930 41870
rect 35534 41858 35586 41870
rect 11330 41806 11342 41858
rect 11394 41806 11406 41858
rect 13458 41806 13470 41858
rect 13522 41806 13534 41858
rect 16930 41806 16942 41858
rect 16994 41806 17006 41858
rect 19170 41806 19182 41858
rect 19234 41806 19246 41858
rect 21410 41806 21422 41858
rect 21474 41806 21486 41858
rect 23202 41806 23214 41858
rect 23266 41806 23278 41858
rect 26450 41806 26462 41858
rect 26514 41806 26526 41858
rect 28578 41806 28590 41858
rect 28642 41806 28654 41858
rect 30482 41806 30494 41858
rect 30546 41806 30558 41858
rect 8878 41794 8930 41806
rect 35534 41794 35586 41806
rect 35982 41858 36034 41870
rect 35982 41794 36034 41806
rect 36430 41858 36482 41870
rect 36430 41794 36482 41806
rect 38670 41858 38722 41870
rect 38670 41794 38722 41806
rect 39118 41858 39170 41870
rect 39118 41794 39170 41806
rect 39566 41858 39618 41870
rect 39566 41794 39618 41806
rect 40014 41858 40066 41870
rect 40014 41794 40066 41806
rect 40462 41858 40514 41870
rect 40462 41794 40514 41806
rect 41470 41858 41522 41870
rect 41470 41794 41522 41806
rect 9886 41746 9938 41758
rect 5506 41694 5518 41746
rect 5570 41743 5582 41746
rect 5842 41743 5854 41746
rect 5570 41697 5854 41743
rect 5570 41694 5582 41697
rect 5842 41694 5854 41697
rect 5906 41743 5918 41746
rect 6066 41743 6078 41746
rect 5906 41697 6078 41743
rect 5906 41694 5918 41697
rect 6066 41694 6078 41697
rect 6130 41743 6142 41746
rect 6290 41743 6302 41746
rect 6130 41697 6302 41743
rect 6130 41694 6142 41697
rect 6290 41694 6302 41697
rect 6354 41694 6366 41746
rect 9886 41682 9938 41694
rect 17950 41746 18002 41758
rect 17950 41682 18002 41694
rect 18174 41746 18226 41758
rect 18174 41682 18226 41694
rect 24446 41746 24498 41758
rect 32062 41746 32114 41758
rect 29922 41694 29934 41746
rect 29986 41694 29998 41746
rect 24446 41682 24498 41694
rect 32062 41682 32114 41694
rect 32286 41746 32338 41758
rect 32286 41682 32338 41694
rect 32510 41746 32562 41758
rect 32510 41682 32562 41694
rect 32622 41746 32674 41758
rect 32622 41682 32674 41694
rect 33630 41746 33682 41758
rect 33630 41682 33682 41694
rect 33966 41746 34018 41758
rect 33966 41682 34018 41694
rect 35086 41746 35138 41758
rect 35970 41694 35982 41746
rect 36034 41743 36046 41746
rect 36754 41743 36766 41746
rect 36034 41697 36766 41743
rect 36034 41694 36046 41697
rect 36754 41694 36766 41697
rect 36818 41694 36830 41746
rect 38882 41694 38894 41746
rect 38946 41743 38958 41746
rect 39666 41743 39678 41746
rect 38946 41697 39678 41743
rect 38946 41694 38958 41697
rect 39666 41694 39678 41697
rect 39730 41694 39742 41746
rect 35086 41682 35138 41694
rect 1344 41578 48608 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 48608 41578
rect 1344 41492 48608 41526
rect 2594 41358 2606 41410
rect 2658 41407 2670 41410
rect 3042 41407 3054 41410
rect 2658 41361 3054 41407
rect 2658 41358 2670 41361
rect 3042 41358 3054 41361
rect 3106 41358 3118 41410
rect 2830 41298 2882 41310
rect 2830 41234 2882 41246
rect 3278 41298 3330 41310
rect 3278 41234 3330 41246
rect 4062 41298 4114 41310
rect 4062 41234 4114 41246
rect 4510 41298 4562 41310
rect 4510 41234 4562 41246
rect 9326 41298 9378 41310
rect 34414 41298 34466 41310
rect 9986 41246 9998 41298
rect 10050 41246 10062 41298
rect 14466 41246 14478 41298
rect 14530 41246 14542 41298
rect 23650 41246 23662 41298
rect 23714 41246 23726 41298
rect 25330 41246 25342 41298
rect 25394 41246 25406 41298
rect 26898 41246 26910 41298
rect 26962 41246 26974 41298
rect 29586 41246 29598 41298
rect 29650 41246 29662 41298
rect 9326 41234 9378 41246
rect 34414 41234 34466 41246
rect 34974 41298 35026 41310
rect 34974 41234 35026 41246
rect 38782 41298 38834 41310
rect 38782 41234 38834 41246
rect 39678 41298 39730 41310
rect 39678 41234 39730 41246
rect 40574 41298 40626 41310
rect 40574 41234 40626 41246
rect 2382 41186 2434 41198
rect 2382 41122 2434 41134
rect 6078 41186 6130 41198
rect 6078 41122 6130 41134
rect 7758 41186 7810 41198
rect 9438 41186 9490 41198
rect 14590 41186 14642 41198
rect 33070 41186 33122 41198
rect 8642 41134 8654 41186
rect 8706 41134 8718 41186
rect 8978 41134 8990 41186
rect 9042 41134 9054 41186
rect 12898 41134 12910 41186
rect 12962 41134 12974 41186
rect 15250 41134 15262 41186
rect 15314 41134 15326 41186
rect 15586 41134 15598 41186
rect 15650 41134 15662 41186
rect 17042 41134 17054 41186
rect 17106 41134 17118 41186
rect 17490 41134 17502 41186
rect 17554 41134 17566 41186
rect 18498 41134 18510 41186
rect 18562 41134 18574 41186
rect 18946 41134 18958 41186
rect 19010 41134 19022 41186
rect 19954 41134 19966 41186
rect 20018 41134 20030 41186
rect 21746 41134 21758 41186
rect 21810 41134 21822 41186
rect 22642 41134 22654 41186
rect 22706 41134 22718 41186
rect 24210 41134 24222 41186
rect 24274 41134 24286 41186
rect 24658 41134 24670 41186
rect 24722 41134 24734 41186
rect 26674 41134 26686 41186
rect 26738 41134 26750 41186
rect 27682 41134 27694 41186
rect 27746 41134 27758 41186
rect 28242 41134 28254 41186
rect 28306 41134 28318 41186
rect 31714 41134 31726 41186
rect 31778 41134 31790 41186
rect 32386 41134 32398 41186
rect 32450 41134 32462 41186
rect 7758 41122 7810 41134
rect 9438 41122 9490 41134
rect 14590 41122 14642 41134
rect 33070 41122 33122 41134
rect 34638 41186 34690 41198
rect 36642 41134 36654 41186
rect 36706 41134 36718 41186
rect 34638 41122 34690 41134
rect 6638 41074 6690 41086
rect 6638 41010 6690 41022
rect 6974 41074 7026 41086
rect 6974 41010 7026 41022
rect 7534 41074 7586 41086
rect 16718 41074 16770 41086
rect 12114 41022 12126 41074
rect 12178 41022 12190 41074
rect 14018 41022 14030 41074
rect 14082 41022 14094 41074
rect 16034 41022 16046 41074
rect 16098 41022 16110 41074
rect 7534 41010 7586 41022
rect 16718 41010 16770 41022
rect 20862 41074 20914 41086
rect 33294 41074 33346 41086
rect 27010 41022 27022 41074
rect 27074 41022 27086 41074
rect 20862 41010 20914 41022
rect 33294 41010 33346 41022
rect 33406 41074 33458 41086
rect 35870 41074 35922 41086
rect 33506 41022 33518 41074
rect 33570 41022 33582 41074
rect 33406 41010 33458 41022
rect 35870 41010 35922 41022
rect 38334 41074 38386 41086
rect 38334 41010 38386 41022
rect 40126 41074 40178 41086
rect 40126 41010 40178 41022
rect 1934 40962 1986 40974
rect 1934 40898 1986 40910
rect 3726 40962 3778 40974
rect 3726 40898 3778 40910
rect 5070 40962 5122 40974
rect 5070 40898 5122 40910
rect 5742 40962 5794 40974
rect 9214 40962 9266 40974
rect 8082 40910 8094 40962
rect 8146 40910 8158 40962
rect 5742 40898 5794 40910
rect 9214 40898 9266 40910
rect 13806 40962 13858 40974
rect 13806 40898 13858 40910
rect 17838 40962 17890 40974
rect 17838 40898 17890 40910
rect 20750 40962 20802 40974
rect 20750 40898 20802 40910
rect 28702 40962 28754 40974
rect 28702 40898 28754 40910
rect 33182 40962 33234 40974
rect 33182 40898 33234 40910
rect 35534 40962 35586 40974
rect 35534 40898 35586 40910
rect 36430 40962 36482 40974
rect 36430 40898 36482 40910
rect 37438 40962 37490 40974
rect 37438 40898 37490 40910
rect 37886 40962 37938 40974
rect 37886 40898 37938 40910
rect 39230 40962 39282 40974
rect 39230 40898 39282 40910
rect 1344 40794 48608 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 48608 40794
rect 1344 40708 48608 40742
rect 2158 40626 2210 40638
rect 2158 40562 2210 40574
rect 3502 40626 3554 40638
rect 3502 40562 3554 40574
rect 5630 40626 5682 40638
rect 5630 40562 5682 40574
rect 6078 40626 6130 40638
rect 6078 40562 6130 40574
rect 9662 40626 9714 40638
rect 18174 40626 18226 40638
rect 9662 40562 9714 40574
rect 9998 40570 10050 40582
rect 3054 40514 3106 40526
rect 3054 40450 3106 40462
rect 6638 40514 6690 40526
rect 6638 40450 6690 40462
rect 7534 40514 7586 40526
rect 7534 40450 7586 40462
rect 8430 40514 8482 40526
rect 8430 40450 8482 40462
rect 9886 40514 9938 40526
rect 18174 40562 18226 40574
rect 19630 40626 19682 40638
rect 31502 40626 31554 40638
rect 23538 40574 23550 40626
rect 23602 40574 23614 40626
rect 19630 40562 19682 40574
rect 31502 40562 31554 40574
rect 34750 40626 34802 40638
rect 34750 40562 34802 40574
rect 35534 40626 35586 40638
rect 35534 40562 35586 40574
rect 35982 40626 36034 40638
rect 35982 40562 36034 40574
rect 37774 40626 37826 40638
rect 37774 40562 37826 40574
rect 38222 40626 38274 40638
rect 38222 40562 38274 40574
rect 9998 40506 10050 40518
rect 48078 40514 48130 40526
rect 22978 40462 22990 40514
rect 23042 40462 23054 40514
rect 24434 40462 24446 40514
rect 24498 40462 24510 40514
rect 26450 40462 26462 40514
rect 26514 40462 26526 40514
rect 29250 40462 29262 40514
rect 29314 40462 29326 40514
rect 30258 40462 30270 40514
rect 30322 40462 30334 40514
rect 9886 40450 9938 40462
rect 48078 40450 48130 40462
rect 3950 40402 4002 40414
rect 3950 40338 4002 40350
rect 4398 40402 4450 40414
rect 4398 40338 4450 40350
rect 6974 40402 7026 40414
rect 6974 40338 7026 40350
rect 7870 40402 7922 40414
rect 17614 40402 17666 40414
rect 10546 40350 10558 40402
rect 10610 40350 10622 40402
rect 11330 40350 11342 40402
rect 11394 40350 11406 40402
rect 14130 40350 14142 40402
rect 14194 40350 14206 40402
rect 14802 40350 14814 40402
rect 14866 40350 14878 40402
rect 7870 40338 7922 40350
rect 17614 40338 17666 40350
rect 18062 40402 18114 40414
rect 18062 40338 18114 40350
rect 18286 40402 18338 40414
rect 19966 40402 20018 40414
rect 19170 40350 19182 40402
rect 19234 40350 19246 40402
rect 18286 40338 18338 40350
rect 19966 40338 20018 40350
rect 20750 40402 20802 40414
rect 32622 40402 32674 40414
rect 21186 40350 21198 40402
rect 21250 40350 21262 40402
rect 22194 40350 22206 40402
rect 22258 40350 22270 40402
rect 22866 40350 22878 40402
rect 22930 40350 22942 40402
rect 24546 40350 24558 40402
rect 24610 40350 24622 40402
rect 25778 40350 25790 40402
rect 25842 40350 25854 40402
rect 29362 40350 29374 40402
rect 29426 40350 29438 40402
rect 30034 40350 30046 40402
rect 30098 40350 30110 40402
rect 30930 40350 30942 40402
rect 30994 40350 31006 40402
rect 20750 40338 20802 40350
rect 32622 40338 32674 40350
rect 33966 40402 34018 40414
rect 33966 40338 34018 40350
rect 34190 40402 34242 40414
rect 34190 40338 34242 40350
rect 35086 40402 35138 40414
rect 35086 40338 35138 40350
rect 36430 40402 36482 40414
rect 36430 40338 36482 40350
rect 39118 40402 39170 40414
rect 39118 40338 39170 40350
rect 39566 40402 39618 40414
rect 39566 40338 39618 40350
rect 2606 40290 2658 40302
rect 2606 40226 2658 40238
rect 4734 40290 4786 40302
rect 4734 40226 4786 40238
rect 5294 40290 5346 40302
rect 18846 40290 18898 40302
rect 32286 40290 32338 40302
rect 13458 40238 13470 40290
rect 13522 40238 13534 40290
rect 16930 40238 16942 40290
rect 16994 40238 17006 40290
rect 28578 40238 28590 40290
rect 28642 40238 28654 40290
rect 5294 40226 5346 40238
rect 18846 40226 18898 40238
rect 32286 40226 32338 40238
rect 36878 40290 36930 40302
rect 36878 40226 36930 40238
rect 37326 40290 37378 40302
rect 37326 40226 37378 40238
rect 38670 40290 38722 40302
rect 38670 40226 38722 40238
rect 8654 40178 8706 40190
rect 3826 40126 3838 40178
rect 3890 40175 3902 40178
rect 4722 40175 4734 40178
rect 3890 40129 4734 40175
rect 3890 40126 3902 40129
rect 4722 40126 4734 40129
rect 4786 40175 4798 40178
rect 5058 40175 5070 40178
rect 4786 40129 5070 40175
rect 4786 40126 4798 40129
rect 5058 40126 5070 40129
rect 5122 40126 5134 40178
rect 8654 40114 8706 40126
rect 8990 40178 9042 40190
rect 8990 40114 9042 40126
rect 31950 40178 32002 40190
rect 31950 40114 32002 40126
rect 32062 40178 32114 40190
rect 32062 40114 32114 40126
rect 32510 40178 32562 40190
rect 32510 40114 32562 40126
rect 33630 40178 33682 40190
rect 33630 40114 33682 40126
rect 1344 40010 48608 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 48608 40010
rect 1344 39924 48608 39958
rect 9102 39842 9154 39854
rect 7074 39790 7086 39842
rect 7138 39839 7150 39842
rect 7634 39839 7646 39842
rect 7138 39793 7646 39839
rect 7138 39790 7150 39793
rect 7634 39790 7646 39793
rect 7698 39790 7710 39842
rect 9102 39778 9154 39790
rect 28702 39842 28754 39854
rect 28702 39778 28754 39790
rect 29598 39842 29650 39854
rect 29598 39778 29650 39790
rect 29822 39842 29874 39854
rect 29822 39778 29874 39790
rect 32510 39842 32562 39854
rect 34850 39790 34862 39842
rect 34914 39839 34926 39842
rect 35186 39839 35198 39842
rect 34914 39793 35198 39839
rect 34914 39790 34926 39793
rect 35186 39790 35198 39793
rect 35250 39790 35262 39842
rect 32510 39778 32562 39790
rect 1822 39730 1874 39742
rect 1822 39666 1874 39678
rect 2382 39730 2434 39742
rect 2382 39666 2434 39678
rect 2830 39730 2882 39742
rect 2830 39666 2882 39678
rect 3614 39730 3666 39742
rect 3614 39666 3666 39678
rect 4510 39730 4562 39742
rect 4510 39666 4562 39678
rect 5630 39730 5682 39742
rect 5630 39666 5682 39678
rect 6190 39730 6242 39742
rect 6190 39666 6242 39678
rect 7086 39730 7138 39742
rect 7086 39666 7138 39678
rect 8094 39730 8146 39742
rect 31166 39730 31218 39742
rect 12898 39678 12910 39730
rect 12962 39678 12974 39730
rect 14466 39678 14478 39730
rect 14530 39678 14542 39730
rect 20850 39678 20862 39730
rect 20914 39678 20926 39730
rect 24546 39678 24558 39730
rect 24610 39678 24622 39730
rect 25106 39678 25118 39730
rect 25170 39678 25182 39730
rect 8094 39666 8146 39678
rect 31166 39666 31218 39678
rect 31390 39730 31442 39742
rect 31390 39666 31442 39678
rect 33070 39730 33122 39742
rect 35534 39730 35586 39742
rect 33730 39678 33742 39730
rect 33794 39678 33806 39730
rect 33070 39666 33122 39678
rect 35534 39666 35586 39678
rect 37886 39730 37938 39742
rect 37886 39666 37938 39678
rect 3278 39618 3330 39630
rect 28590 39618 28642 39630
rect 30270 39618 30322 39630
rect 32846 39618 32898 39630
rect 38334 39618 38386 39630
rect 10098 39566 10110 39618
rect 10162 39566 10174 39618
rect 17266 39566 17278 39618
rect 17330 39566 17342 39618
rect 17938 39566 17950 39618
rect 18002 39566 18014 39618
rect 21634 39566 21646 39618
rect 21698 39566 21710 39618
rect 27906 39566 27918 39618
rect 27970 39566 27982 39618
rect 30146 39566 30158 39618
rect 30210 39566 30222 39618
rect 31714 39566 31726 39618
rect 31778 39566 31790 39618
rect 33618 39566 33630 39618
rect 33682 39566 33694 39618
rect 3278 39554 3330 39566
rect 28590 39554 28642 39566
rect 30270 39554 30322 39566
rect 32846 39554 32898 39566
rect 38334 39554 38386 39566
rect 38782 39618 38834 39630
rect 38782 39554 38834 39566
rect 7982 39506 8034 39518
rect 7982 39442 8034 39454
rect 8878 39506 8930 39518
rect 13582 39506 13634 39518
rect 10770 39454 10782 39506
rect 10834 39454 10846 39506
rect 8878 39442 8930 39454
rect 13582 39442 13634 39454
rect 13918 39506 13970 39518
rect 33966 39506 34018 39518
rect 16594 39454 16606 39506
rect 16658 39454 16670 39506
rect 18722 39454 18734 39506
rect 18786 39454 18798 39506
rect 22418 39454 22430 39506
rect 22482 39454 22494 39506
rect 27234 39454 27246 39506
rect 27298 39454 27310 39506
rect 13918 39442 13970 39454
rect 33966 39442 34018 39454
rect 34638 39506 34690 39518
rect 34638 39442 34690 39454
rect 35086 39506 35138 39518
rect 35086 39442 35138 39454
rect 4174 39394 4226 39406
rect 4174 39330 4226 39342
rect 5070 39394 5122 39406
rect 5070 39330 5122 39342
rect 6526 39394 6578 39406
rect 6526 39330 6578 39342
rect 7422 39394 7474 39406
rect 7422 39330 7474 39342
rect 8206 39394 8258 39406
rect 13806 39394 13858 39406
rect 9426 39342 9438 39394
rect 9490 39342 9502 39394
rect 8206 39330 8258 39342
rect 13806 39330 13858 39342
rect 28702 39394 28754 39406
rect 28702 39330 28754 39342
rect 30382 39394 30434 39406
rect 30382 39330 30434 39342
rect 30494 39394 30546 39406
rect 30494 39330 30546 39342
rect 34526 39394 34578 39406
rect 34526 39330 34578 39342
rect 35982 39394 36034 39406
rect 35982 39330 36034 39342
rect 36430 39394 36482 39406
rect 36430 39330 36482 39342
rect 37438 39394 37490 39406
rect 37438 39330 37490 39342
rect 1344 39226 48608 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 48608 39226
rect 1344 39140 48608 39174
rect 3726 39058 3778 39070
rect 3726 38994 3778 39006
rect 5070 39058 5122 39070
rect 5070 38994 5122 39006
rect 5854 39058 5906 39070
rect 5854 38994 5906 39006
rect 7758 39058 7810 39070
rect 7758 38994 7810 39006
rect 9102 39058 9154 39070
rect 9102 38994 9154 39006
rect 10222 39058 10274 39070
rect 33518 39058 33570 39070
rect 11778 39006 11790 39058
rect 11842 39006 11854 39058
rect 10222 38994 10274 39006
rect 33518 38994 33570 39006
rect 34414 39058 34466 39070
rect 34414 38994 34466 39006
rect 35758 39058 35810 39070
rect 35758 38994 35810 39006
rect 36206 39058 36258 39070
rect 36206 38994 36258 39006
rect 36654 39058 36706 39070
rect 36654 38994 36706 39006
rect 37102 39058 37154 39070
rect 37102 38994 37154 39006
rect 1822 38946 1874 38958
rect 1822 38882 1874 38894
rect 6414 38946 6466 38958
rect 21422 38946 21474 38958
rect 29262 38946 29314 38958
rect 29710 38946 29762 38958
rect 14802 38894 14814 38946
rect 14866 38894 14878 38946
rect 20402 38894 20414 38946
rect 20466 38894 20478 38946
rect 27794 38894 27806 38946
rect 27858 38894 27870 38946
rect 29474 38894 29486 38946
rect 29538 38894 29550 38946
rect 6414 38882 6466 38894
rect 21422 38882 21474 38894
rect 29262 38882 29314 38894
rect 29710 38882 29762 38894
rect 31278 38946 31330 38958
rect 31278 38882 31330 38894
rect 32174 38946 32226 38958
rect 32174 38882 32226 38894
rect 32846 38946 32898 38958
rect 32846 38882 32898 38894
rect 37550 38946 37602 38958
rect 37550 38882 37602 38894
rect 4174 38834 4226 38846
rect 4174 38770 4226 38782
rect 10222 38834 10274 38846
rect 10222 38770 10274 38782
rect 10334 38834 10386 38846
rect 10334 38770 10386 38782
rect 10558 38834 10610 38846
rect 19742 38834 19794 38846
rect 30046 38834 30098 38846
rect 12898 38782 12910 38834
rect 12962 38782 12974 38834
rect 14130 38782 14142 38834
rect 14194 38782 14206 38834
rect 18274 38782 18286 38834
rect 18338 38782 18350 38834
rect 19170 38782 19182 38834
rect 19234 38782 19246 38834
rect 20514 38782 20526 38834
rect 20578 38782 20590 38834
rect 21074 38782 21086 38834
rect 21138 38782 21150 38834
rect 21970 38782 21982 38834
rect 22034 38782 22046 38834
rect 28466 38782 28478 38834
rect 28530 38782 28542 38834
rect 10558 38770 10610 38782
rect 19742 38770 19794 38782
rect 30046 38770 30098 38782
rect 30158 38834 30210 38846
rect 30158 38770 30210 38782
rect 31726 38834 31778 38846
rect 31726 38770 31778 38782
rect 32398 38834 32450 38846
rect 32398 38770 32450 38782
rect 33966 38834 34018 38846
rect 33966 38770 34018 38782
rect 35310 38834 35362 38846
rect 35310 38770 35362 38782
rect 4622 38722 4674 38734
rect 4622 38658 4674 38670
rect 5518 38722 5570 38734
rect 5518 38658 5570 38670
rect 6750 38722 6802 38734
rect 6750 38658 6802 38670
rect 7310 38722 7362 38734
rect 7310 38658 7362 38670
rect 8094 38722 8146 38734
rect 8094 38658 8146 38670
rect 8542 38722 8594 38734
rect 8542 38658 8594 38670
rect 11230 38722 11282 38734
rect 11230 38658 11282 38670
rect 11454 38722 11506 38734
rect 13358 38722 13410 38734
rect 17614 38722 17666 38734
rect 31950 38722 32002 38734
rect 13010 38670 13022 38722
rect 13074 38670 13086 38722
rect 16930 38670 16942 38722
rect 16994 38670 17006 38722
rect 22754 38670 22766 38722
rect 22818 38670 22830 38722
rect 24882 38670 24894 38722
rect 24946 38670 24958 38722
rect 25666 38670 25678 38722
rect 25730 38670 25742 38722
rect 29138 38670 29150 38722
rect 29202 38670 29214 38722
rect 11454 38658 11506 38670
rect 13358 38658 13410 38670
rect 17614 38658 17666 38670
rect 31950 38658 32002 38670
rect 34862 38722 34914 38734
rect 34862 38658 34914 38670
rect 30718 38610 30770 38622
rect 17602 38558 17614 38610
rect 17666 38607 17678 38610
rect 17938 38607 17950 38610
rect 17666 38561 17950 38607
rect 17666 38558 17678 38561
rect 17938 38558 17950 38561
rect 18002 38558 18014 38610
rect 30718 38546 30770 38558
rect 31054 38610 31106 38622
rect 32498 38558 32510 38610
rect 32562 38607 32574 38610
rect 32722 38607 32734 38610
rect 32562 38561 32734 38607
rect 32562 38558 32574 38561
rect 32722 38558 32734 38561
rect 32786 38558 32798 38610
rect 33506 38558 33518 38610
rect 33570 38607 33582 38610
rect 34178 38607 34190 38610
rect 33570 38561 34190 38607
rect 33570 38558 33582 38561
rect 34178 38558 34190 38561
rect 34242 38558 34254 38610
rect 31054 38546 31106 38558
rect 1344 38442 48608 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 48608 38442
rect 1344 38356 48608 38390
rect 12350 38274 12402 38286
rect 6850 38222 6862 38274
rect 6914 38271 6926 38274
rect 7522 38271 7534 38274
rect 6914 38225 7534 38271
rect 6914 38222 6926 38225
rect 7522 38222 7534 38225
rect 7586 38222 7598 38274
rect 7746 38222 7758 38274
rect 7810 38271 7822 38274
rect 8194 38271 8206 38274
rect 7810 38225 8206 38271
rect 7810 38222 7822 38225
rect 8194 38222 8206 38225
rect 8258 38222 8270 38274
rect 12350 38210 12402 38222
rect 30158 38274 30210 38286
rect 30158 38210 30210 38222
rect 32174 38274 32226 38286
rect 32386 38222 32398 38274
rect 32450 38271 32462 38274
rect 33170 38271 33182 38274
rect 32450 38225 33182 38271
rect 32450 38222 32462 38225
rect 33170 38222 33182 38225
rect 33234 38271 33246 38274
rect 34066 38271 34078 38274
rect 33234 38225 34078 38271
rect 33234 38222 33246 38225
rect 34066 38222 34078 38225
rect 34130 38222 34142 38274
rect 35746 38222 35758 38274
rect 35810 38271 35822 38274
rect 36642 38271 36654 38274
rect 35810 38225 36654 38271
rect 35810 38222 35822 38225
rect 36642 38222 36654 38225
rect 36706 38222 36718 38274
rect 32174 38210 32226 38222
rect 4062 38162 4114 38174
rect 4062 38098 4114 38110
rect 4622 38162 4674 38174
rect 4622 38098 4674 38110
rect 5854 38162 5906 38174
rect 5854 38098 5906 38110
rect 6638 38162 6690 38174
rect 6638 38098 6690 38110
rect 9886 38162 9938 38174
rect 33070 38162 33122 38174
rect 17378 38110 17390 38162
rect 17442 38110 17454 38162
rect 20850 38110 20862 38162
rect 20914 38110 20926 38162
rect 24546 38110 24558 38162
rect 24610 38110 24622 38162
rect 28018 38110 28030 38162
rect 28082 38110 28094 38162
rect 9886 38098 9938 38110
rect 33070 38098 33122 38110
rect 36206 38162 36258 38174
rect 36206 38098 36258 38110
rect 10670 38050 10722 38062
rect 12574 38050 12626 38062
rect 12114 37998 12126 38050
rect 12178 37998 12190 38050
rect 10670 37986 10722 37998
rect 12574 37986 12626 37998
rect 12798 38050 12850 38062
rect 12798 37986 12850 37998
rect 14030 38050 14082 38062
rect 29822 38050 29874 38062
rect 14578 37998 14590 38050
rect 14642 37998 14654 38050
rect 17938 37998 17950 38050
rect 18002 37998 18014 38050
rect 21634 37998 21646 38050
rect 21698 37998 21710 38050
rect 25218 37998 25230 38050
rect 25282 37998 25294 38050
rect 14030 37986 14082 37998
rect 29822 37986 29874 37998
rect 30942 38050 30994 38062
rect 30942 37986 30994 37998
rect 32622 38050 32674 38062
rect 32622 37986 32674 37998
rect 35758 38050 35810 38062
rect 35758 37986 35810 37998
rect 5070 37938 5122 37950
rect 5070 37874 5122 37886
rect 7534 37938 7586 37950
rect 7534 37874 7586 37886
rect 7982 37938 8034 37950
rect 7982 37874 8034 37886
rect 8430 37938 8482 37950
rect 8430 37874 8482 37886
rect 10334 37938 10386 37950
rect 10334 37874 10386 37886
rect 13694 37938 13746 37950
rect 28590 37938 28642 37950
rect 15250 37886 15262 37938
rect 15314 37886 15326 37938
rect 18722 37886 18734 37938
rect 18786 37886 18798 37938
rect 22418 37886 22430 37938
rect 22482 37886 22494 37938
rect 25890 37886 25902 37938
rect 25954 37886 25966 37938
rect 13694 37874 13746 37886
rect 28590 37874 28642 37886
rect 29598 37938 29650 37950
rect 29598 37874 29650 37886
rect 30718 37938 30770 37950
rect 30718 37874 30770 37886
rect 31278 37938 31330 37950
rect 31278 37874 31330 37886
rect 31950 37938 32002 37950
rect 31950 37874 32002 37886
rect 33966 37938 34018 37950
rect 33966 37874 34018 37886
rect 6302 37826 6354 37838
rect 6302 37762 6354 37774
rect 7198 37826 7250 37838
rect 7198 37762 7250 37774
rect 8990 37826 9042 37838
rect 8990 37762 9042 37774
rect 9326 37826 9378 37838
rect 11566 37826 11618 37838
rect 11218 37774 11230 37826
rect 11282 37774 11294 37826
rect 9326 37762 9378 37774
rect 11566 37762 11618 37774
rect 12238 37826 12290 37838
rect 12238 37762 12290 37774
rect 13806 37826 13858 37838
rect 13806 37762 13858 37774
rect 28702 37826 28754 37838
rect 28702 37762 28754 37774
rect 28926 37826 28978 37838
rect 28926 37762 28978 37774
rect 30830 37826 30882 37838
rect 30830 37762 30882 37774
rect 32062 37826 32114 37838
rect 32062 37762 32114 37774
rect 33518 37826 33570 37838
rect 33518 37762 33570 37774
rect 34414 37826 34466 37838
rect 34414 37762 34466 37774
rect 34862 37826 34914 37838
rect 34862 37762 34914 37774
rect 35310 37826 35362 37838
rect 35310 37762 35362 37774
rect 36654 37826 36706 37838
rect 36654 37762 36706 37774
rect 48078 37826 48130 37838
rect 48078 37762 48130 37774
rect 1344 37658 48608 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 48608 37658
rect 1344 37572 48608 37606
rect 5966 37490 6018 37502
rect 5966 37426 6018 37438
rect 6302 37490 6354 37502
rect 6302 37426 6354 37438
rect 7758 37490 7810 37502
rect 7758 37426 7810 37438
rect 8654 37490 8706 37502
rect 8654 37426 8706 37438
rect 9998 37490 10050 37502
rect 9998 37426 10050 37438
rect 11454 37490 11506 37502
rect 11454 37426 11506 37438
rect 12238 37490 12290 37502
rect 31278 37490 31330 37502
rect 18050 37438 18062 37490
rect 18114 37438 18126 37490
rect 12238 37426 12290 37438
rect 31278 37426 31330 37438
rect 32734 37490 32786 37502
rect 32734 37426 32786 37438
rect 34862 37490 34914 37502
rect 34862 37426 34914 37438
rect 1822 37378 1874 37390
rect 28702 37378 28754 37390
rect 30158 37378 30210 37390
rect 16146 37326 16158 37378
rect 16210 37326 16222 37378
rect 18386 37326 18398 37378
rect 18450 37326 18462 37378
rect 18610 37326 18622 37378
rect 18674 37326 18686 37378
rect 23874 37326 23886 37378
rect 23938 37326 23950 37378
rect 25890 37326 25902 37378
rect 25954 37326 25966 37378
rect 27234 37326 27246 37378
rect 27298 37326 27310 37378
rect 29250 37326 29262 37378
rect 29314 37326 29326 37378
rect 1822 37314 1874 37326
rect 28702 37314 28754 37326
rect 30158 37314 30210 37326
rect 30382 37378 30434 37390
rect 30382 37314 30434 37326
rect 33966 37378 34018 37390
rect 33966 37314 34018 37326
rect 6862 37266 6914 37278
rect 6862 37202 6914 37214
rect 11118 37266 11170 37278
rect 11118 37202 11170 37214
rect 13470 37266 13522 37278
rect 28590 37266 28642 37278
rect 16818 37214 16830 37266
rect 16882 37214 16894 37266
rect 18946 37214 18958 37266
rect 19010 37214 19022 37266
rect 22306 37214 22318 37266
rect 22370 37214 22382 37266
rect 27010 37214 27022 37266
rect 27074 37214 27086 37266
rect 13470 37202 13522 37214
rect 28590 37202 28642 37214
rect 28814 37266 28866 37278
rect 28814 37202 28866 37214
rect 29710 37266 29762 37278
rect 29710 37202 29762 37214
rect 30942 37266 30994 37278
rect 30942 37202 30994 37214
rect 33518 37266 33570 37278
rect 33518 37202 33570 37214
rect 5518 37154 5570 37166
rect 5518 37090 5570 37102
rect 7198 37154 7250 37166
rect 7198 37090 7250 37102
rect 8206 37154 8258 37166
rect 8206 37090 8258 37102
rect 8990 37154 9042 37166
rect 8990 37090 9042 37102
rect 10446 37154 10498 37166
rect 25678 37154 25730 37166
rect 12338 37102 12350 37154
rect 12402 37102 12414 37154
rect 14018 37102 14030 37154
rect 14082 37102 14094 37154
rect 19506 37102 19518 37154
rect 19570 37102 19582 37154
rect 21634 37102 21646 37154
rect 21698 37102 21710 37154
rect 23986 37102 23998 37154
rect 24050 37102 24062 37154
rect 10446 37090 10498 37102
rect 25678 37090 25730 37102
rect 29934 37154 29986 37166
rect 29934 37090 29986 37102
rect 31726 37154 31778 37166
rect 31726 37090 31778 37102
rect 32174 37154 32226 37166
rect 32174 37090 32226 37102
rect 34414 37154 34466 37166
rect 34414 37090 34466 37102
rect 35310 37154 35362 37166
rect 35310 37090 35362 37102
rect 35758 37154 35810 37166
rect 35758 37090 35810 37102
rect 10558 37042 10610 37054
rect 10558 36978 10610 36990
rect 12014 37042 12066 37054
rect 12014 36978 12066 36990
rect 12910 37042 12962 37054
rect 12910 36978 12962 36990
rect 13246 37042 13298 37054
rect 13246 36978 13298 36990
rect 23102 37042 23154 37054
rect 35298 36990 35310 37042
rect 35362 37039 35374 37042
rect 35634 37039 35646 37042
rect 35362 36993 35646 37039
rect 35362 36990 35374 36993
rect 35634 36990 35646 36993
rect 35698 36990 35710 37042
rect 23102 36978 23154 36990
rect 1344 36874 48608 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 48608 36874
rect 1344 36788 48608 36822
rect 6962 36654 6974 36706
rect 7026 36703 7038 36706
rect 7634 36703 7646 36706
rect 7026 36657 7646 36703
rect 7026 36654 7038 36657
rect 7634 36654 7646 36657
rect 7698 36654 7710 36706
rect 8978 36654 8990 36706
rect 9042 36703 9054 36706
rect 9314 36703 9326 36706
rect 9042 36657 9326 36703
rect 9042 36654 9054 36657
rect 9314 36654 9326 36657
rect 9378 36654 9390 36706
rect 26114 36654 26126 36706
rect 26178 36654 26190 36706
rect 30370 36654 30382 36706
rect 30434 36703 30446 36706
rect 31378 36703 31390 36706
rect 30434 36657 31390 36703
rect 30434 36654 30446 36657
rect 31378 36654 31390 36657
rect 31442 36654 31454 36706
rect 34626 36654 34638 36706
rect 34690 36703 34702 36706
rect 34850 36703 34862 36706
rect 34690 36657 34862 36703
rect 34690 36654 34702 36657
rect 34850 36654 34862 36657
rect 34914 36654 34926 36706
rect 6302 36594 6354 36606
rect 6302 36530 6354 36542
rect 7646 36594 7698 36606
rect 7646 36530 7698 36542
rect 8430 36594 8482 36606
rect 8430 36530 8482 36542
rect 8878 36594 8930 36606
rect 8878 36530 8930 36542
rect 10222 36594 10274 36606
rect 10222 36530 10274 36542
rect 10670 36594 10722 36606
rect 27470 36594 27522 36606
rect 15250 36542 15262 36594
rect 15314 36542 15326 36594
rect 17378 36542 17390 36594
rect 17442 36542 17454 36594
rect 17938 36542 17950 36594
rect 18002 36542 18014 36594
rect 21634 36542 21646 36594
rect 21698 36542 21710 36594
rect 23762 36542 23774 36594
rect 23826 36542 23838 36594
rect 26002 36542 26014 36594
rect 26066 36542 26078 36594
rect 10670 36530 10722 36542
rect 27470 36530 27522 36542
rect 31390 36594 31442 36606
rect 31390 36530 31442 36542
rect 32734 36594 32786 36606
rect 32734 36530 32786 36542
rect 34078 36594 34130 36606
rect 34078 36530 34130 36542
rect 34862 36594 34914 36606
rect 34862 36530 34914 36542
rect 14030 36482 14082 36494
rect 27134 36482 27186 36494
rect 14578 36430 14590 36482
rect 14642 36430 14654 36482
rect 20066 36430 20078 36482
rect 20130 36430 20142 36482
rect 20738 36430 20750 36482
rect 20802 36430 20814 36482
rect 24434 36430 24446 36482
rect 24498 36430 24510 36482
rect 25330 36430 25342 36482
rect 25394 36430 25406 36482
rect 14030 36418 14082 36430
rect 27134 36418 27186 36430
rect 27246 36482 27298 36494
rect 27246 36418 27298 36430
rect 28590 36482 28642 36494
rect 30382 36482 30434 36494
rect 29586 36430 29598 36482
rect 29650 36430 29662 36482
rect 28590 36418 28642 36430
rect 30382 36418 30434 36430
rect 9326 36370 9378 36382
rect 9326 36306 9378 36318
rect 11230 36370 11282 36382
rect 11230 36306 11282 36318
rect 11678 36370 11730 36382
rect 11678 36306 11730 36318
rect 12910 36370 12962 36382
rect 12910 36306 12962 36318
rect 13694 36370 13746 36382
rect 13694 36306 13746 36318
rect 13806 36370 13858 36382
rect 13806 36306 13858 36318
rect 26798 36370 26850 36382
rect 26798 36306 26850 36318
rect 27694 36370 27746 36382
rect 27694 36306 27746 36318
rect 28254 36370 28306 36382
rect 28254 36306 28306 36318
rect 28814 36370 28866 36382
rect 28814 36306 28866 36318
rect 29934 36370 29986 36382
rect 29934 36306 29986 36318
rect 31726 36370 31778 36382
rect 31726 36306 31778 36318
rect 6750 36258 6802 36270
rect 6750 36194 6802 36206
rect 7086 36258 7138 36270
rect 7086 36194 7138 36206
rect 7982 36258 8034 36270
rect 7982 36194 8034 36206
rect 9774 36258 9826 36270
rect 9774 36194 9826 36206
rect 12014 36258 12066 36270
rect 12014 36194 12066 36206
rect 12574 36258 12626 36270
rect 12574 36194 12626 36206
rect 27806 36258 27858 36270
rect 27806 36194 27858 36206
rect 28366 36258 28418 36270
rect 28366 36194 28418 36206
rect 29822 36258 29874 36270
rect 29822 36194 29874 36206
rect 30830 36258 30882 36270
rect 30830 36194 30882 36206
rect 32174 36258 32226 36270
rect 32174 36194 32226 36206
rect 33070 36258 33122 36270
rect 33070 36194 33122 36206
rect 33630 36258 33682 36270
rect 33630 36194 33682 36206
rect 34414 36258 34466 36270
rect 34414 36194 34466 36206
rect 48078 36258 48130 36270
rect 48078 36194 48130 36206
rect 1344 36090 48608 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 48608 36090
rect 1344 36004 48608 36038
rect 8094 35922 8146 35934
rect 8094 35858 8146 35870
rect 8990 35922 9042 35934
rect 8990 35858 9042 35870
rect 10782 35922 10834 35934
rect 10782 35858 10834 35870
rect 13582 35922 13634 35934
rect 13582 35858 13634 35870
rect 14478 35922 14530 35934
rect 14478 35858 14530 35870
rect 15486 35922 15538 35934
rect 18846 35922 18898 35934
rect 16594 35870 16606 35922
rect 16658 35870 16670 35922
rect 15486 35858 15538 35870
rect 18846 35858 18898 35870
rect 22878 35922 22930 35934
rect 22878 35858 22930 35870
rect 26462 35922 26514 35934
rect 29150 35922 29202 35934
rect 27122 35870 27134 35922
rect 27186 35870 27198 35922
rect 26462 35858 26514 35870
rect 29150 35858 29202 35870
rect 30606 35922 30658 35934
rect 30606 35858 30658 35870
rect 31950 35922 32002 35934
rect 31950 35858 32002 35870
rect 32846 35922 32898 35934
rect 32846 35858 32898 35870
rect 33518 35922 33570 35934
rect 33518 35858 33570 35870
rect 1822 35810 1874 35822
rect 1822 35746 1874 35758
rect 12574 35810 12626 35822
rect 12574 35746 12626 35758
rect 14142 35810 14194 35822
rect 14142 35746 14194 35758
rect 17726 35810 17778 35822
rect 28254 35810 28306 35822
rect 20066 35758 20078 35810
rect 20130 35758 20142 35810
rect 24210 35758 24222 35810
rect 24274 35758 24286 35810
rect 25890 35758 25902 35810
rect 25954 35758 25966 35810
rect 17726 35746 17778 35758
rect 28254 35746 28306 35758
rect 28590 35810 28642 35822
rect 28590 35746 28642 35758
rect 29262 35810 29314 35822
rect 29262 35746 29314 35758
rect 32398 35810 32450 35822
rect 32398 35746 32450 35758
rect 8654 35698 8706 35710
rect 8654 35634 8706 35646
rect 13246 35698 13298 35710
rect 13246 35634 13298 35646
rect 15038 35698 15090 35710
rect 15038 35634 15090 35646
rect 15374 35698 15426 35710
rect 15374 35634 15426 35646
rect 15598 35698 15650 35710
rect 15598 35634 15650 35646
rect 16158 35698 16210 35710
rect 18174 35698 18226 35710
rect 26350 35698 26402 35710
rect 16370 35646 16382 35698
rect 16434 35646 16446 35698
rect 16930 35646 16942 35698
rect 16994 35646 17006 35698
rect 19282 35646 19294 35698
rect 19346 35646 19358 35698
rect 22866 35646 22878 35698
rect 22930 35646 22942 35698
rect 23314 35646 23326 35698
rect 23378 35646 23390 35698
rect 23986 35646 23998 35698
rect 24050 35646 24062 35698
rect 25666 35646 25678 35698
rect 25730 35646 25742 35698
rect 16158 35634 16210 35646
rect 18174 35634 18226 35646
rect 26350 35634 26402 35646
rect 26574 35698 26626 35710
rect 26574 35634 26626 35646
rect 31502 35698 31554 35710
rect 31502 35634 31554 35646
rect 7310 35586 7362 35598
rect 7310 35522 7362 35534
rect 7758 35586 7810 35598
rect 7758 35522 7810 35534
rect 9886 35586 9938 35598
rect 9886 35522 9938 35534
rect 10222 35586 10274 35598
rect 10222 35522 10274 35534
rect 11230 35586 11282 35598
rect 11230 35522 11282 35534
rect 11678 35586 11730 35598
rect 11678 35522 11730 35534
rect 12014 35586 12066 35598
rect 24782 35586 24834 35598
rect 22194 35534 22206 35586
rect 22258 35534 22270 35586
rect 12014 35522 12066 35534
rect 24782 35522 24834 35534
rect 24894 35586 24946 35598
rect 24894 35522 24946 35534
rect 27470 35586 27522 35598
rect 27470 35522 27522 35534
rect 27694 35586 27746 35598
rect 27694 35522 27746 35534
rect 29710 35586 29762 35598
rect 29710 35522 29762 35534
rect 30158 35586 30210 35598
rect 30158 35522 30210 35534
rect 31166 35586 31218 35598
rect 31166 35522 31218 35534
rect 12686 35474 12738 35486
rect 12686 35410 12738 35422
rect 16606 35474 16658 35486
rect 16606 35410 16658 35422
rect 17950 35474 18002 35486
rect 17950 35410 18002 35422
rect 18398 35474 18450 35486
rect 18398 35410 18450 35422
rect 26126 35474 26178 35486
rect 30370 35422 30382 35474
rect 30434 35471 30446 35474
rect 31826 35471 31838 35474
rect 30434 35425 31838 35471
rect 30434 35422 30446 35425
rect 31826 35422 31838 35425
rect 31890 35422 31902 35474
rect 26126 35410 26178 35422
rect 1344 35306 48608 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 48608 35306
rect 1344 35220 48608 35254
rect 16494 35138 16546 35150
rect 9314 35086 9326 35138
rect 9378 35135 9390 35138
rect 9762 35135 9774 35138
rect 9378 35089 9774 35135
rect 9378 35086 9390 35089
rect 9762 35086 9774 35089
rect 9826 35086 9838 35138
rect 11666 35086 11678 35138
rect 11730 35135 11742 35138
rect 12002 35135 12014 35138
rect 11730 35089 12014 35135
rect 11730 35086 11742 35089
rect 12002 35086 12014 35089
rect 12066 35086 12078 35138
rect 16494 35074 16546 35086
rect 25454 35138 25506 35150
rect 25454 35074 25506 35086
rect 25678 35138 25730 35150
rect 25678 35074 25730 35086
rect 27918 35138 27970 35150
rect 30146 35086 30158 35138
rect 30210 35135 30222 35138
rect 32722 35135 32734 35138
rect 30210 35089 32734 35135
rect 30210 35086 30222 35089
rect 32722 35086 32734 35089
rect 32786 35086 32798 35138
rect 27918 35074 27970 35086
rect 8878 35026 8930 35038
rect 8878 34962 8930 34974
rect 9326 35026 9378 35038
rect 9326 34962 9378 34974
rect 9774 35026 9826 35038
rect 9774 34962 9826 34974
rect 10334 35026 10386 35038
rect 10334 34962 10386 34974
rect 12014 35026 12066 35038
rect 29934 35026 29986 35038
rect 14914 34974 14926 35026
rect 14978 34974 14990 35026
rect 15698 34974 15710 35026
rect 15762 34974 15774 35026
rect 17938 34974 17950 35026
rect 18002 34974 18014 35026
rect 21634 34974 21646 35026
rect 21698 34974 21710 35026
rect 12014 34962 12066 34974
rect 29934 34962 29986 34974
rect 30942 35026 30994 35038
rect 30942 34962 30994 34974
rect 31390 35026 31442 35038
rect 31390 34962 31442 34974
rect 31726 35026 31778 35038
rect 31726 34962 31778 34974
rect 11230 34914 11282 34926
rect 11230 34850 11282 34862
rect 11566 34914 11618 34926
rect 16942 34914 16994 34926
rect 15810 34862 15822 34914
rect 15874 34862 15886 34914
rect 11566 34850 11618 34862
rect 16942 34850 16994 34862
rect 17166 34914 17218 34926
rect 17166 34850 17218 34862
rect 17390 34914 17442 34926
rect 25230 34914 25282 34926
rect 20738 34862 20750 34914
rect 20802 34862 20814 34914
rect 24434 34862 24446 34914
rect 24498 34862 24510 34914
rect 17390 34850 17442 34862
rect 25230 34850 25282 34862
rect 25790 34914 25842 34926
rect 25790 34850 25842 34862
rect 26798 34914 26850 34926
rect 26798 34850 26850 34862
rect 28590 34914 28642 34926
rect 28590 34850 28642 34862
rect 30494 34914 30546 34926
rect 30494 34850 30546 34862
rect 13806 34802 13858 34814
rect 13806 34738 13858 34750
rect 14142 34802 14194 34814
rect 14142 34738 14194 34750
rect 14702 34802 14754 34814
rect 14702 34738 14754 34750
rect 15598 34802 15650 34814
rect 15598 34738 15650 34750
rect 16046 34802 16098 34814
rect 27022 34802 27074 34814
rect 20066 34750 20078 34802
rect 20130 34750 20142 34802
rect 23762 34750 23774 34802
rect 23826 34750 23838 34802
rect 16046 34738 16098 34750
rect 27022 34738 27074 34750
rect 27694 34802 27746 34814
rect 27694 34738 27746 34750
rect 10670 34690 10722 34702
rect 10670 34626 10722 34638
rect 12574 34690 12626 34702
rect 12574 34626 12626 34638
rect 13022 34690 13074 34702
rect 13022 34626 13074 34638
rect 14926 34690 14978 34702
rect 14926 34626 14978 34638
rect 25342 34690 25394 34702
rect 27806 34690 27858 34702
rect 26450 34638 26462 34690
rect 26514 34638 26526 34690
rect 25342 34626 25394 34638
rect 27806 34626 27858 34638
rect 28478 34690 28530 34702
rect 28478 34626 28530 34638
rect 29598 34690 29650 34702
rect 29598 34626 29650 34638
rect 32174 34690 32226 34702
rect 32174 34626 32226 34638
rect 32734 34690 32786 34702
rect 32734 34626 32786 34638
rect 48078 34690 48130 34702
rect 48078 34626 48130 34638
rect 1344 34522 48608 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 48608 34522
rect 1344 34436 48608 34470
rect 9774 34354 9826 34366
rect 9774 34290 9826 34302
rect 10222 34354 10274 34366
rect 10222 34290 10274 34302
rect 11006 34354 11058 34366
rect 11006 34290 11058 34302
rect 11566 34354 11618 34366
rect 11566 34290 11618 34302
rect 12014 34354 12066 34366
rect 12014 34290 12066 34302
rect 12462 34354 12514 34366
rect 12462 34290 12514 34302
rect 12910 34354 12962 34366
rect 12910 34290 12962 34302
rect 13694 34354 13746 34366
rect 13694 34290 13746 34302
rect 15038 34354 15090 34366
rect 24670 34354 24722 34366
rect 15922 34302 15934 34354
rect 15986 34302 15998 34354
rect 15038 34290 15090 34302
rect 24670 34290 24722 34302
rect 26574 34354 26626 34366
rect 26574 34290 26626 34302
rect 27470 34354 27522 34366
rect 27470 34290 27522 34302
rect 28030 34354 28082 34366
rect 28030 34290 28082 34302
rect 28478 34354 28530 34366
rect 28478 34290 28530 34302
rect 29822 34354 29874 34366
rect 29822 34290 29874 34302
rect 30382 34354 30434 34366
rect 30382 34290 30434 34302
rect 30718 34354 30770 34366
rect 30718 34290 30770 34302
rect 31166 34354 31218 34366
rect 31166 34290 31218 34302
rect 16494 34242 16546 34254
rect 16494 34178 16546 34190
rect 25678 34242 25730 34254
rect 25678 34178 25730 34190
rect 26014 34242 26066 34254
rect 26014 34178 26066 34190
rect 26910 34242 26962 34254
rect 26910 34178 26962 34190
rect 27582 34242 27634 34254
rect 27582 34178 27634 34190
rect 13246 34130 13298 34142
rect 13246 34066 13298 34078
rect 14702 34130 14754 34142
rect 14702 34066 14754 34078
rect 15598 34130 15650 34142
rect 17054 34130 17106 34142
rect 16706 34078 16718 34130
rect 16770 34078 16782 34130
rect 15598 34066 15650 34078
rect 17054 34066 17106 34078
rect 18062 34130 18114 34142
rect 18062 34066 18114 34078
rect 18286 34130 18338 34142
rect 24446 34130 24498 34142
rect 29374 34130 29426 34142
rect 19170 34078 19182 34130
rect 19234 34078 19246 34130
rect 23090 34078 23102 34130
rect 23154 34078 23166 34130
rect 24210 34078 24222 34130
rect 24274 34078 24286 34130
rect 24882 34078 24894 34130
rect 24946 34078 24958 34130
rect 27906 34078 27918 34130
rect 27970 34078 27982 34130
rect 18286 34066 18338 34078
rect 24446 34066 24498 34078
rect 10558 34018 10610 34030
rect 10558 33954 10610 33966
rect 14142 34018 14194 34030
rect 16594 33966 16606 34018
rect 16658 33966 16670 34018
rect 19842 33966 19854 34018
rect 19906 33966 19918 34018
rect 21970 33966 21982 34018
rect 22034 33966 22046 34018
rect 23426 33966 23438 34018
rect 23490 33966 23502 34018
rect 24770 33966 24782 34018
rect 24834 33966 24846 34018
rect 14142 33954 14194 33966
rect 17726 33906 17778 33918
rect 17726 33842 17778 33854
rect 17838 33906 17890 33918
rect 17838 33842 17890 33854
rect 18398 33906 18450 33918
rect 23538 33854 23550 33906
rect 23602 33854 23614 33906
rect 27921 33903 27967 34078
rect 29374 34066 29426 34078
rect 28926 34018 28978 34030
rect 28926 33954 28978 33966
rect 28914 33903 28926 33906
rect 27921 33857 28926 33903
rect 28914 33854 28926 33857
rect 28978 33903 28990 33906
rect 30146 33903 30158 33906
rect 28978 33857 30158 33903
rect 28978 33854 28990 33857
rect 30146 33854 30158 33857
rect 30210 33854 30222 33906
rect 18398 33842 18450 33854
rect 1344 33738 48608 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 48608 33738
rect 1344 33652 48608 33686
rect 23774 33570 23826 33582
rect 3490 33518 3502 33570
rect 3554 33567 3566 33570
rect 4162 33567 4174 33570
rect 3554 33521 4174 33567
rect 3554 33518 3566 33521
rect 4162 33518 4174 33521
rect 4226 33518 4238 33570
rect 13682 33518 13694 33570
rect 13746 33567 13758 33570
rect 15026 33567 15038 33570
rect 13746 33521 15038 33567
rect 13746 33518 13758 33521
rect 15026 33518 15038 33521
rect 15090 33518 15102 33570
rect 19394 33518 19406 33570
rect 19458 33518 19470 33570
rect 23774 33506 23826 33518
rect 24558 33570 24610 33582
rect 27682 33518 27694 33570
rect 27746 33567 27758 33570
rect 27906 33567 27918 33570
rect 27746 33521 27918 33567
rect 27746 33518 27758 33521
rect 27906 33518 27918 33521
rect 27970 33518 27982 33570
rect 24558 33506 24610 33518
rect 3838 33458 3890 33470
rect 3838 33394 3890 33406
rect 11006 33458 11058 33470
rect 11006 33394 11058 33406
rect 11678 33458 11730 33470
rect 11678 33394 11730 33406
rect 12126 33458 12178 33470
rect 12126 33394 12178 33406
rect 12574 33458 12626 33470
rect 12574 33394 12626 33406
rect 14142 33458 14194 33470
rect 14142 33394 14194 33406
rect 15486 33458 15538 33470
rect 15486 33394 15538 33406
rect 15822 33458 15874 33470
rect 15822 33394 15874 33406
rect 18622 33458 18674 33470
rect 20862 33458 20914 33470
rect 26350 33458 26402 33470
rect 20066 33406 20078 33458
rect 20130 33406 20142 33458
rect 21858 33406 21870 33458
rect 21922 33406 21934 33458
rect 24770 33406 24782 33458
rect 24834 33406 24846 33458
rect 18622 33394 18674 33406
rect 20862 33394 20914 33406
rect 26350 33394 26402 33406
rect 26910 33458 26962 33470
rect 26910 33394 26962 33406
rect 27470 33458 27522 33470
rect 27470 33394 27522 33406
rect 27918 33458 27970 33470
rect 27918 33394 27970 33406
rect 28814 33458 28866 33470
rect 28814 33394 28866 33406
rect 29486 33458 29538 33470
rect 29486 33394 29538 33406
rect 4734 33346 4786 33358
rect 4734 33282 4786 33294
rect 15038 33346 15090 33358
rect 22654 33346 22706 33358
rect 17378 33294 17390 33346
rect 17442 33294 17454 33346
rect 19730 33294 19742 33346
rect 19794 33294 19806 33346
rect 21970 33294 21982 33346
rect 22034 33294 22046 33346
rect 15038 33282 15090 33294
rect 22654 33282 22706 33294
rect 23326 33346 23378 33358
rect 23326 33282 23378 33294
rect 23550 33346 23602 33358
rect 23550 33282 23602 33294
rect 23886 33346 23938 33358
rect 25666 33294 25678 33346
rect 25730 33294 25742 33346
rect 23886 33282 23938 33294
rect 4398 33234 4450 33246
rect 4398 33170 4450 33182
rect 14590 33234 14642 33246
rect 14590 33170 14642 33182
rect 23214 33234 23266 33246
rect 23214 33170 23266 33182
rect 24782 33234 24834 33246
rect 24782 33170 24834 33182
rect 25454 33234 25506 33246
rect 25454 33170 25506 33182
rect 28366 33234 28418 33246
rect 28366 33170 28418 33182
rect 1822 33122 1874 33134
rect 1822 33058 1874 33070
rect 13022 33122 13074 33134
rect 13022 33058 13074 33070
rect 13582 33122 13634 33134
rect 16718 33122 16770 33134
rect 16370 33070 16382 33122
rect 16434 33070 16446 33122
rect 13582 33058 13634 33070
rect 16718 33058 16770 33070
rect 17614 33122 17666 33134
rect 17614 33058 17666 33070
rect 18286 33122 18338 33134
rect 18286 33058 18338 33070
rect 18510 33122 18562 33134
rect 18510 33058 18562 33070
rect 18734 33122 18786 33134
rect 18734 33058 18786 33070
rect 26462 33122 26514 33134
rect 26462 33058 26514 33070
rect 1344 32954 48608 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 48608 32954
rect 1344 32868 48608 32902
rect 12574 32786 12626 32798
rect 12574 32722 12626 32734
rect 14926 32786 14978 32798
rect 14926 32722 14978 32734
rect 16158 32786 16210 32798
rect 16158 32722 16210 32734
rect 16830 32786 16882 32798
rect 16830 32722 16882 32734
rect 17054 32786 17106 32798
rect 22206 32786 22258 32798
rect 18834 32734 18846 32786
rect 18898 32734 18910 32786
rect 17054 32722 17106 32734
rect 22206 32722 22258 32734
rect 22318 32786 22370 32798
rect 22318 32722 22370 32734
rect 25678 32786 25730 32798
rect 25678 32722 25730 32734
rect 26014 32786 26066 32798
rect 26014 32722 26066 32734
rect 27022 32786 27074 32798
rect 27022 32722 27074 32734
rect 27470 32786 27522 32798
rect 27470 32722 27522 32734
rect 27918 32786 27970 32798
rect 27918 32722 27970 32734
rect 28366 32786 28418 32798
rect 28366 32722 28418 32734
rect 13582 32674 13634 32686
rect 13582 32610 13634 32622
rect 16718 32674 16770 32686
rect 16718 32610 16770 32622
rect 19406 32674 19458 32686
rect 19406 32610 19458 32622
rect 21086 32674 21138 32686
rect 21086 32610 21138 32622
rect 22430 32674 22482 32686
rect 22430 32610 22482 32622
rect 22542 32674 22594 32686
rect 22542 32610 22594 32622
rect 23550 32674 23602 32686
rect 23550 32610 23602 32622
rect 23998 32674 24050 32686
rect 23998 32610 24050 32622
rect 24558 32674 24610 32686
rect 24558 32610 24610 32622
rect 24894 32674 24946 32686
rect 24894 32610 24946 32622
rect 48078 32674 48130 32686
rect 48078 32610 48130 32622
rect 15374 32562 15426 32574
rect 15374 32498 15426 32510
rect 19742 32562 19794 32574
rect 20974 32562 21026 32574
rect 20178 32510 20190 32562
rect 20242 32510 20254 32562
rect 22978 32510 22990 32562
rect 23042 32510 23054 32562
rect 23762 32510 23774 32562
rect 23826 32510 23838 32562
rect 19742 32498 19794 32510
rect 20974 32498 21026 32510
rect 12238 32450 12290 32462
rect 12238 32386 12290 32398
rect 13134 32450 13186 32462
rect 13134 32386 13186 32398
rect 14030 32450 14082 32462
rect 14030 32386 14082 32398
rect 14478 32450 14530 32462
rect 14478 32386 14530 32398
rect 15710 32450 15762 32462
rect 15710 32386 15762 32398
rect 17726 32450 17778 32462
rect 17726 32386 17778 32398
rect 18286 32450 18338 32462
rect 18286 32386 18338 32398
rect 23662 32450 23714 32462
rect 23662 32386 23714 32398
rect 26574 32450 26626 32462
rect 26574 32386 26626 32398
rect 18510 32338 18562 32350
rect 18510 32274 18562 32286
rect 19518 32338 19570 32350
rect 19518 32274 19570 32286
rect 19966 32338 20018 32350
rect 19966 32274 20018 32286
rect 20750 32338 20802 32350
rect 20750 32274 20802 32286
rect 21310 32338 21362 32350
rect 21310 32274 21362 32286
rect 21534 32338 21586 32350
rect 21534 32274 21586 32286
rect 1344 32170 48608 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 48608 32170
rect 1344 32084 48608 32118
rect 14254 31890 14306 31902
rect 14254 31826 14306 31838
rect 15598 31890 15650 31902
rect 15598 31826 15650 31838
rect 21870 31890 21922 31902
rect 21870 31826 21922 31838
rect 22878 31890 22930 31902
rect 22878 31826 22930 31838
rect 24670 31890 24722 31902
rect 24670 31826 24722 31838
rect 25230 31890 25282 31902
rect 25230 31826 25282 31838
rect 25678 31890 25730 31902
rect 25678 31826 25730 31838
rect 27022 31890 27074 31902
rect 27022 31826 27074 31838
rect 16382 31778 16434 31790
rect 19182 31778 19234 31790
rect 18498 31726 18510 31778
rect 18562 31726 18574 31778
rect 16382 31714 16434 31726
rect 19182 31714 19234 31726
rect 20190 31778 20242 31790
rect 20190 31714 20242 31726
rect 20302 31778 20354 31790
rect 20302 31714 20354 31726
rect 21646 31778 21698 31790
rect 21646 31714 21698 31726
rect 22654 31778 22706 31790
rect 22654 31714 22706 31726
rect 26574 31778 26626 31790
rect 26574 31714 26626 31726
rect 16046 31666 16098 31678
rect 16046 31602 16098 31614
rect 18286 31666 18338 31678
rect 18286 31602 18338 31614
rect 20414 31666 20466 31678
rect 20414 31602 20466 31614
rect 23214 31666 23266 31678
rect 23214 31602 23266 31614
rect 24110 31666 24162 31678
rect 24110 31602 24162 31614
rect 14702 31554 14754 31566
rect 14702 31490 14754 31502
rect 15150 31554 15202 31566
rect 15150 31490 15202 31502
rect 16942 31554 16994 31566
rect 16942 31490 16994 31502
rect 17278 31554 17330 31566
rect 17278 31490 17330 31502
rect 17838 31554 17890 31566
rect 17838 31490 17890 31502
rect 19518 31554 19570 31566
rect 22990 31554 23042 31566
rect 20850 31502 20862 31554
rect 20914 31502 20926 31554
rect 22194 31502 22206 31554
rect 22258 31502 22270 31554
rect 19518 31490 19570 31502
rect 22990 31490 23042 31502
rect 23774 31554 23826 31566
rect 23774 31490 23826 31502
rect 26126 31554 26178 31566
rect 26126 31490 26178 31502
rect 48078 31554 48130 31566
rect 48078 31490 48130 31502
rect 1344 31386 48608 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 48608 31386
rect 1344 31300 48608 31334
rect 14814 31218 14866 31230
rect 14814 31154 14866 31166
rect 16606 31218 16658 31230
rect 16606 31154 16658 31166
rect 17054 31218 17106 31230
rect 17054 31154 17106 31166
rect 18510 31218 18562 31230
rect 18510 31154 18562 31166
rect 19742 31218 19794 31230
rect 23550 31218 23602 31230
rect 23314 31166 23326 31218
rect 23378 31166 23390 31218
rect 19742 31154 19794 31166
rect 19070 31106 19122 31118
rect 19070 31042 19122 31054
rect 19518 31106 19570 31118
rect 19518 31042 19570 31054
rect 22990 31106 23042 31118
rect 22990 31042 23042 31054
rect 15598 30994 15650 31006
rect 15598 30930 15650 30942
rect 18174 30994 18226 31006
rect 18174 30930 18226 30942
rect 21870 30994 21922 31006
rect 22754 30942 22766 30994
rect 22818 30942 22830 30994
rect 21870 30930 21922 30942
rect 16158 30882 16210 30894
rect 16158 30818 16210 30830
rect 17726 30882 17778 30894
rect 17726 30818 17778 30830
rect 22094 30882 22146 30894
rect 22094 30818 22146 30830
rect 19854 30770 19906 30782
rect 16146 30718 16158 30770
rect 16210 30767 16222 30770
rect 16482 30767 16494 30770
rect 16210 30721 16494 30767
rect 16210 30718 16222 30721
rect 16482 30718 16494 30721
rect 16546 30767 16558 30770
rect 16706 30767 16718 30770
rect 16546 30721 16718 30767
rect 16546 30718 16558 30721
rect 16706 30718 16718 30721
rect 16770 30718 16782 30770
rect 19854 30706 19906 30718
rect 20414 30770 20466 30782
rect 20414 30706 20466 30718
rect 20526 30770 20578 30782
rect 20526 30706 20578 30718
rect 20750 30770 20802 30782
rect 20750 30706 20802 30718
rect 20862 30770 20914 30782
rect 20862 30706 20914 30718
rect 21534 30770 21586 30782
rect 23329 30770 23375 31166
rect 23550 31154 23602 31166
rect 24894 31218 24946 31230
rect 24894 31154 24946 31166
rect 25678 31218 25730 31230
rect 25678 31154 25730 31166
rect 23998 31106 24050 31118
rect 23998 31042 24050 31054
rect 24446 30882 24498 30894
rect 24446 30818 24498 30830
rect 26126 30882 26178 30894
rect 26126 30818 26178 30830
rect 23314 30718 23326 30770
rect 23378 30718 23390 30770
rect 21534 30706 21586 30718
rect 1344 30602 48608 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 48608 30602
rect 1344 30516 48608 30550
rect 22194 30382 22206 30434
rect 22258 30431 22270 30434
rect 22754 30431 22766 30434
rect 22258 30385 22766 30431
rect 22258 30382 22270 30385
rect 22754 30382 22766 30385
rect 22818 30431 22830 30434
rect 23426 30431 23438 30434
rect 22818 30385 23438 30431
rect 22818 30382 22830 30385
rect 23426 30382 23438 30385
rect 23490 30382 23502 30434
rect 17278 30322 17330 30334
rect 17278 30258 17330 30270
rect 17838 30322 17890 30334
rect 17838 30258 17890 30270
rect 19630 30322 19682 30334
rect 19630 30258 19682 30270
rect 23438 30322 23490 30334
rect 23438 30258 23490 30270
rect 24334 30322 24386 30334
rect 24334 30258 24386 30270
rect 16158 30210 16210 30222
rect 16158 30146 16210 30158
rect 18286 30210 18338 30222
rect 18286 30146 18338 30158
rect 19182 30210 19234 30222
rect 19182 30146 19234 30158
rect 20078 30210 20130 30222
rect 20078 30146 20130 30158
rect 23886 30210 23938 30222
rect 23886 30146 23938 30158
rect 25118 30210 25170 30222
rect 25118 30146 25170 30158
rect 20862 30098 20914 30110
rect 20862 30034 20914 30046
rect 21982 30098 22034 30110
rect 21982 30034 22034 30046
rect 1822 29986 1874 29998
rect 1822 29922 1874 29934
rect 18734 29986 18786 29998
rect 18734 29922 18786 29934
rect 20526 29986 20578 29998
rect 20526 29922 20578 29934
rect 21646 29986 21698 29998
rect 21646 29922 21698 29934
rect 22430 29986 22482 29998
rect 22430 29922 22482 29934
rect 22878 29986 22930 29998
rect 22878 29922 22930 29934
rect 24782 29986 24834 29998
rect 24782 29922 24834 29934
rect 1344 29818 48608 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 48608 29818
rect 1344 29732 48608 29766
rect 19182 29650 19234 29662
rect 19182 29586 19234 29598
rect 19742 29650 19794 29662
rect 19742 29586 19794 29598
rect 20750 29650 20802 29662
rect 20750 29586 20802 29598
rect 21198 29650 21250 29662
rect 21198 29586 21250 29598
rect 21982 29650 22034 29662
rect 21982 29586 22034 29598
rect 22542 29650 22594 29662
rect 22542 29586 22594 29598
rect 22990 29650 23042 29662
rect 22990 29586 23042 29598
rect 23438 29650 23490 29662
rect 23438 29586 23490 29598
rect 23886 29650 23938 29662
rect 23886 29586 23938 29598
rect 48078 29538 48130 29550
rect 48078 29474 48130 29486
rect 20302 29314 20354 29326
rect 20302 29250 20354 29262
rect 21646 29314 21698 29326
rect 21646 29250 21698 29262
rect 20290 29150 20302 29202
rect 20354 29199 20366 29202
rect 20626 29199 20638 29202
rect 20354 29153 20638 29199
rect 20354 29150 20366 29153
rect 20626 29150 20638 29153
rect 20690 29150 20702 29202
rect 21970 29150 21982 29202
rect 22034 29199 22046 29202
rect 22530 29199 22542 29202
rect 22034 29153 22542 29199
rect 22034 29150 22046 29153
rect 22530 29150 22542 29153
rect 22594 29150 22606 29202
rect 1344 29034 48608 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 48608 29034
rect 1344 28948 48608 28982
rect 21982 28754 22034 28766
rect 21982 28690 22034 28702
rect 22542 28754 22594 28766
rect 22542 28690 22594 28702
rect 22990 28754 23042 28766
rect 22990 28690 23042 28702
rect 1822 28418 1874 28430
rect 1822 28354 1874 28366
rect 1344 28250 48608 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 48608 28250
rect 1344 28164 48608 28198
rect 1344 27466 48608 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 48608 27466
rect 1344 27380 48608 27414
rect 1822 26850 1874 26862
rect 1822 26786 1874 26798
rect 48078 26850 48130 26862
rect 48078 26786 48130 26798
rect 1344 26682 48608 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 48608 26682
rect 1344 26596 48608 26630
rect 1344 25898 48608 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 48608 25898
rect 1344 25812 48608 25846
rect 1344 25114 48608 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 48608 25114
rect 1344 25028 48608 25062
rect 1822 24834 1874 24846
rect 1822 24770 1874 24782
rect 1344 24330 48608 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 48608 24330
rect 1344 24244 48608 24278
rect 48078 23714 48130 23726
rect 48078 23650 48130 23662
rect 1344 23546 48608 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 48608 23546
rect 1344 23460 48608 23494
rect 3502 23378 3554 23390
rect 3502 23314 3554 23326
rect 3042 23102 3054 23154
rect 3106 23102 3118 23154
rect 2034 22990 2046 23042
rect 2098 22990 2110 23042
rect 1344 22762 48608 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 48608 22762
rect 1344 22676 48608 22710
rect 48078 22146 48130 22158
rect 48078 22082 48130 22094
rect 1344 21978 48608 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 48608 21978
rect 1344 21892 48608 21926
rect 1822 21698 1874 21710
rect 1822 21634 1874 21646
rect 1344 21194 48608 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 48608 21194
rect 1344 21108 48608 21142
rect 1344 20410 48608 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 48608 20410
rect 1344 20324 48608 20358
rect 1344 19626 48608 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 48608 19626
rect 1344 19540 48608 19574
rect 1822 19010 1874 19022
rect 1822 18946 1874 18958
rect 1344 18842 48608 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 48608 18842
rect 1344 18756 48608 18790
rect 48078 18562 48130 18574
rect 48078 18498 48130 18510
rect 1344 18058 48608 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 48608 18058
rect 1344 17972 48608 18006
rect 1822 17554 1874 17566
rect 1822 17490 1874 17502
rect 48078 17442 48130 17454
rect 48078 17378 48130 17390
rect 1344 17274 48608 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 48608 17274
rect 1344 17188 48608 17222
rect 1344 16490 48608 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 48608 16490
rect 1344 16404 48608 16438
rect 1822 15874 1874 15886
rect 1822 15810 1874 15822
rect 1344 15706 48608 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 48608 15706
rect 1344 15620 48608 15654
rect 1344 14922 48608 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 48608 14922
rect 1344 14836 48608 14870
rect 1822 14306 1874 14318
rect 1822 14242 1874 14254
rect 1344 14138 48608 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 48608 14138
rect 1344 14052 48608 14086
rect 1344 13354 48608 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 48608 13354
rect 1344 13268 48608 13302
rect 48078 12850 48130 12862
rect 48078 12786 48130 12798
rect 1344 12570 48608 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 48608 12570
rect 1344 12484 48608 12518
rect 48078 12290 48130 12302
rect 48078 12226 48130 12238
rect 1344 11786 48608 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 48608 11786
rect 1344 11700 48608 11734
rect 1344 11002 48608 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 48608 11002
rect 1344 10916 48608 10950
rect 1822 10722 1874 10734
rect 1822 10658 1874 10670
rect 1344 10218 48608 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 48608 10218
rect 1344 10132 48608 10166
rect 9102 9714 9154 9726
rect 9102 9650 9154 9662
rect 8766 9602 8818 9614
rect 8766 9538 8818 9550
rect 9550 9602 9602 9614
rect 9550 9538 9602 9550
rect 48078 9602 48130 9614
rect 48078 9538 48130 9550
rect 1344 9434 48608 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 48608 9434
rect 1344 9348 48608 9382
rect 1822 9154 1874 9166
rect 1822 9090 1874 9102
rect 1344 8650 48608 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 48608 8650
rect 1344 8564 48608 8598
rect 48078 8034 48130 8046
rect 48078 7970 48130 7982
rect 1344 7866 48608 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 48608 7866
rect 1344 7780 48608 7814
rect 1822 7586 1874 7598
rect 1822 7522 1874 7534
rect 1344 7082 48608 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 48608 7082
rect 1344 6996 48608 7030
rect 48078 6466 48130 6478
rect 48078 6402 48130 6414
rect 1344 6298 48608 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 48608 6298
rect 1344 6212 48608 6246
rect 1344 5514 48608 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 48608 5514
rect 1344 5428 48608 5462
rect 1344 4730 48608 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 48608 4730
rect 1344 4644 48608 4678
rect 1822 4450 1874 4462
rect 1822 4386 1874 4398
rect 2494 4450 2546 4462
rect 2494 4386 2546 4398
rect 48078 4450 48130 4462
rect 48078 4386 48130 4398
rect 47518 4226 47570 4238
rect 47518 4162 47570 4174
rect 1344 3946 48608 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 48608 3946
rect 1344 3860 48608 3894
rect 4286 3666 4338 3678
rect 4286 3602 4338 3614
rect 2146 3502 2158 3554
rect 2210 3502 2222 3554
rect 3042 3502 3054 3554
rect 3106 3502 3118 3554
rect 11902 3442 11954 3454
rect 11902 3378 11954 3390
rect 12350 3442 12402 3454
rect 12350 3378 12402 3390
rect 18622 3442 18674 3454
rect 18622 3378 18674 3390
rect 19070 3442 19122 3454
rect 19070 3378 19122 3390
rect 36430 3442 36482 3454
rect 36430 3378 36482 3390
rect 37550 3442 37602 3454
rect 37550 3378 37602 3390
rect 48078 3442 48130 3454
rect 48078 3378 48130 3390
rect 3614 3330 3666 3342
rect 3614 3266 3666 3278
rect 5742 3330 5794 3342
rect 5742 3266 5794 3278
rect 9662 3330 9714 3342
rect 9662 3266 9714 3278
rect 12686 3330 12738 3342
rect 12686 3266 12738 3278
rect 14366 3330 14418 3342
rect 14366 3266 14418 3278
rect 15710 3330 15762 3342
rect 15710 3266 15762 3278
rect 17726 3330 17778 3342
rect 17726 3266 17778 3278
rect 19406 3330 19458 3342
rect 19406 3266 19458 3278
rect 21422 3330 21474 3342
rect 21422 3266 21474 3278
rect 23102 3330 23154 3342
rect 23102 3266 23154 3278
rect 26462 3330 26514 3342
rect 26462 3266 26514 3278
rect 29262 3330 29314 3342
rect 29262 3266 29314 3278
rect 31838 3330 31890 3342
rect 31838 3266 31890 3278
rect 35198 3330 35250 3342
rect 35198 3266 35250 3278
rect 37214 3330 37266 3342
rect 37214 3266 37266 3278
rect 38558 3330 38610 3342
rect 38558 3266 38610 3278
rect 41022 3330 41074 3342
rect 41022 3266 41074 3278
rect 42590 3330 42642 3342
rect 42590 3266 42642 3278
rect 43934 3330 43986 3342
rect 43934 3266 43986 3278
rect 45950 3330 46002 3342
rect 45950 3266 46002 3278
rect 47182 3330 47234 3342
rect 47182 3266 47234 3278
rect 47742 3330 47794 3342
rect 47742 3266 47794 3278
rect 1344 3162 48608 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 48608 3162
rect 1344 3076 48608 3110
rect 40338 1822 40350 1874
rect 40402 1871 40414 1874
rect 41010 1871 41022 1874
rect 40402 1825 41022 1871
rect 40402 1822 40414 1825
rect 41010 1822 41022 1825
rect 41074 1822 41086 1874
rect 8754 1710 8766 1762
rect 8818 1759 8830 1762
rect 9650 1759 9662 1762
rect 8818 1713 9662 1759
rect 8818 1710 8830 1713
rect 9650 1710 9662 1713
rect 9714 1710 9726 1762
rect 20850 1710 20862 1762
rect 20914 1759 20926 1762
rect 21410 1759 21422 1762
rect 20914 1713 21422 1759
rect 20914 1710 20926 1713
rect 21410 1710 21422 1713
rect 21474 1710 21486 1762
<< via1 >>
rect 25566 48974 25618 49026
rect 26462 48974 26514 49026
rect 22990 48750 23042 48802
rect 27022 48750 27074 48802
rect 23662 47742 23714 47794
rect 23998 47742 24050 47794
rect 27022 47742 27074 47794
rect 13918 47406 13970 47458
rect 15486 47406 15538 47458
rect 16718 47406 16770 47458
rect 14702 47182 14754 47234
rect 16046 47182 16098 47234
rect 8318 46958 8370 47010
rect 8542 46958 8594 47010
rect 32286 46734 32338 46786
rect 33406 46734 33458 46786
rect 27694 46510 27746 46562
rect 29822 46510 29874 46562
rect 31950 46510 32002 46562
rect 2046 46398 2098 46450
rect 2718 46398 2770 46450
rect 8878 46398 8930 46450
rect 9438 46398 9490 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 28366 46062 28418 46114
rect 4062 45950 4114 46002
rect 5854 45950 5906 46002
rect 7198 45950 7250 46002
rect 9774 45950 9826 46002
rect 11902 45950 11954 46002
rect 17726 45950 17778 46002
rect 19854 45950 19906 46002
rect 22206 45950 22258 46002
rect 24334 45950 24386 46002
rect 25790 45950 25842 46002
rect 26350 45950 26402 46002
rect 33406 45950 33458 46002
rect 35646 45950 35698 46002
rect 38446 45950 38498 46002
rect 38894 45950 38946 46002
rect 39342 45950 39394 46002
rect 1822 45838 1874 45890
rect 4846 45838 4898 45890
rect 13582 45838 13634 45890
rect 20638 45838 20690 45890
rect 21534 45838 21586 45890
rect 26014 45838 26066 45890
rect 27806 45838 27858 45890
rect 34190 45838 34242 45890
rect 36094 45838 36146 45890
rect 41806 45838 41858 45890
rect 2158 45726 2210 45778
rect 2718 45726 2770 45778
rect 7646 45726 7698 45778
rect 8878 45726 8930 45778
rect 10334 45726 10386 45778
rect 11006 45726 11058 45778
rect 11566 45726 11618 45778
rect 12462 45726 12514 45778
rect 15374 45726 15426 45778
rect 27358 45726 27410 45778
rect 27470 45726 27522 45778
rect 27582 45726 27634 45778
rect 28478 45726 28530 45778
rect 30158 45726 30210 45778
rect 31502 45726 31554 45778
rect 32062 45726 32114 45778
rect 37886 45726 37938 45778
rect 39902 45726 39954 45778
rect 41358 45726 41410 45778
rect 43262 45726 43314 45778
rect 48078 45726 48130 45778
rect 6190 45614 6242 45666
rect 6638 45614 6690 45666
rect 8206 45614 8258 45666
rect 11790 45614 11842 45666
rect 12798 45614 12850 45666
rect 16718 45614 16770 45666
rect 27694 45614 27746 45666
rect 29262 45614 29314 45666
rect 29598 45614 29650 45666
rect 31166 45614 31218 45666
rect 37102 45614 37154 45666
rect 40910 45614 40962 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 1822 45278 1874 45330
rect 2494 45278 2546 45330
rect 3166 45278 3218 45330
rect 4622 45278 4674 45330
rect 5070 45278 5122 45330
rect 5966 45278 6018 45330
rect 8206 45278 8258 45330
rect 8542 45278 8594 45330
rect 9102 45278 9154 45330
rect 10670 45278 10722 45330
rect 12238 45278 12290 45330
rect 31502 45278 31554 45330
rect 32062 45278 32114 45330
rect 32398 45278 32450 45330
rect 36206 45278 36258 45330
rect 37102 45278 37154 45330
rect 38446 45278 38498 45330
rect 39342 45278 39394 45330
rect 39790 45278 39842 45330
rect 40686 45278 40738 45330
rect 11118 45166 11170 45218
rect 11454 45166 11506 45218
rect 13470 45166 13522 45218
rect 18622 45166 18674 45218
rect 22990 45166 23042 45218
rect 26014 45166 26066 45218
rect 28030 45166 28082 45218
rect 28926 45166 28978 45218
rect 29262 45166 29314 45218
rect 30382 45166 30434 45218
rect 34862 45166 34914 45218
rect 6750 45054 6802 45106
rect 13246 45054 13298 45106
rect 14030 45054 14082 45106
rect 17726 45054 17778 45106
rect 19518 45054 19570 45106
rect 23102 45054 23154 45106
rect 23774 45054 23826 45106
rect 24446 45054 24498 45106
rect 25790 45054 25842 45106
rect 26574 45054 26626 45106
rect 28142 45054 28194 45106
rect 28366 45054 28418 45106
rect 29374 45054 29426 45106
rect 30046 45054 30098 45106
rect 33630 45054 33682 45106
rect 4174 44942 4226 44994
rect 5518 44942 5570 44994
rect 6302 44942 6354 44994
rect 7310 44942 7362 44994
rect 7758 44942 7810 44994
rect 9774 44942 9826 44994
rect 10222 44942 10274 44994
rect 12910 44942 12962 44994
rect 14814 44942 14866 44994
rect 16942 44942 16994 44994
rect 20302 44942 20354 44994
rect 22430 44942 22482 44994
rect 24894 44942 24946 44994
rect 27582 44942 27634 44994
rect 29038 44942 29090 44994
rect 31054 44942 31106 44994
rect 32846 44942 32898 44994
rect 33966 44942 34018 44994
rect 34414 44942 34466 44994
rect 35310 44942 35362 44994
rect 35758 44942 35810 44994
rect 36654 44942 36706 44994
rect 37550 44942 37602 44994
rect 37998 44942 38050 44994
rect 38894 44942 38946 44994
rect 40238 44942 40290 44994
rect 12014 44830 12066 44882
rect 12350 44830 12402 44882
rect 24558 44830 24610 44882
rect 26910 44830 26962 44882
rect 30046 44830 30098 44882
rect 30942 44830 30994 44882
rect 31950 44830 32002 44882
rect 32846 44830 32898 44882
rect 36990 44830 37042 44882
rect 37998 44830 38050 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 11454 44494 11506 44546
rect 11790 44494 11842 44546
rect 28702 44494 28754 44546
rect 33966 44494 34018 44546
rect 34638 44494 34690 44546
rect 3726 44382 3778 44434
rect 4174 44382 4226 44434
rect 5070 44382 5122 44434
rect 6750 44382 6802 44434
rect 7198 44382 7250 44434
rect 8094 44382 8146 44434
rect 9774 44382 9826 44434
rect 11230 44382 11282 44434
rect 15262 44382 15314 44434
rect 17390 44382 17442 44434
rect 18734 44382 18786 44434
rect 20862 44382 20914 44434
rect 22430 44382 22482 44434
rect 24558 44382 24610 44434
rect 25902 44382 25954 44434
rect 28030 44382 28082 44434
rect 31166 44382 31218 44434
rect 33070 44382 33122 44434
rect 33966 44382 34018 44434
rect 37438 44382 37490 44434
rect 38334 44382 38386 44434
rect 39678 44382 39730 44434
rect 3054 44270 3106 44322
rect 4622 44270 4674 44322
rect 10446 44270 10498 44322
rect 12350 44270 12402 44322
rect 12910 44270 12962 44322
rect 14030 44270 14082 44322
rect 14478 44270 14530 44322
rect 17950 44270 18002 44322
rect 21646 44270 21698 44322
rect 25230 44270 25282 44322
rect 29822 44270 29874 44322
rect 30718 44270 30770 44322
rect 31054 44270 31106 44322
rect 31838 44270 31890 44322
rect 38782 44270 38834 44322
rect 2158 44158 2210 44210
rect 5854 44158 5906 44210
rect 10670 44158 10722 44210
rect 12574 44158 12626 44210
rect 13694 44158 13746 44210
rect 13806 44158 13858 44210
rect 28702 44158 28754 44210
rect 28814 44158 28866 44210
rect 32174 44158 32226 44210
rect 35310 44158 35362 44210
rect 6190 44046 6242 44098
rect 7646 44046 7698 44098
rect 8430 44046 8482 44098
rect 8990 44046 9042 44098
rect 9438 44046 9490 44098
rect 12686 44046 12738 44098
rect 29598 44046 29650 44098
rect 29710 44046 29762 44098
rect 30046 44046 30098 44098
rect 31278 44046 31330 44098
rect 32734 44046 32786 44098
rect 33518 44046 33570 44098
rect 34526 44046 34578 44098
rect 34974 44046 35026 44098
rect 35758 44046 35810 44098
rect 36206 44046 36258 44098
rect 36654 44046 36706 44098
rect 37886 44046 37938 44098
rect 39230 44046 39282 44098
rect 40126 44046 40178 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 1934 43710 1986 43762
rect 10670 43710 10722 43762
rect 11678 43710 11730 43762
rect 18958 43710 19010 43762
rect 31054 43710 31106 43762
rect 31726 43710 31778 43762
rect 37102 43710 37154 43762
rect 38894 43710 38946 43762
rect 40686 43710 40738 43762
rect 47742 43710 47794 43762
rect 3726 43598 3778 43650
rect 4958 43598 5010 43650
rect 8206 43598 8258 43650
rect 9886 43598 9938 43650
rect 11454 43598 11506 43650
rect 11790 43598 11842 43650
rect 14814 43598 14866 43650
rect 17950 43598 18002 43650
rect 18398 43598 18450 43650
rect 27806 43598 27858 43650
rect 31838 43598 31890 43650
rect 32062 43598 32114 43650
rect 33966 43598 34018 43650
rect 4174 43486 4226 43538
rect 6750 43486 6802 43538
rect 10446 43486 10498 43538
rect 11230 43486 11282 43538
rect 13022 43486 13074 43538
rect 13470 43486 13522 43538
rect 14030 43486 14082 43538
rect 18622 43486 18674 43538
rect 19630 43486 19682 43538
rect 23326 43486 23378 43538
rect 24110 43486 24162 43538
rect 24558 43486 24610 43538
rect 28478 43486 28530 43538
rect 29486 43486 29538 43538
rect 29710 43486 29762 43538
rect 29822 43486 29874 43538
rect 30046 43486 30098 43538
rect 30718 43486 30770 43538
rect 30830 43486 30882 43538
rect 30942 43486 30994 43538
rect 31278 43486 31330 43538
rect 32398 43486 32450 43538
rect 37998 43486 38050 43538
rect 48078 43486 48130 43538
rect 2382 43374 2434 43426
rect 2830 43374 2882 43426
rect 3166 43374 3218 43426
rect 4622 43374 4674 43426
rect 5518 43374 5570 43426
rect 5966 43374 6018 43426
rect 6302 43374 6354 43426
rect 7310 43374 7362 43426
rect 7758 43374 7810 43426
rect 8654 43374 8706 43426
rect 9102 43374 9154 43426
rect 12686 43374 12738 43426
rect 16942 43374 16994 43426
rect 20414 43374 20466 43426
rect 22542 43374 22594 43426
rect 23662 43374 23714 43426
rect 25678 43374 25730 43426
rect 29038 43374 29090 43426
rect 32734 43374 32786 43426
rect 33518 43374 33570 43426
rect 34414 43374 34466 43426
rect 34862 43374 34914 43426
rect 35310 43374 35362 43426
rect 35758 43374 35810 43426
rect 36206 43374 36258 43426
rect 36654 43374 36706 43426
rect 37550 43374 37602 43426
rect 38446 43374 38498 43426
rect 39342 43374 39394 43426
rect 39790 43374 39842 43426
rect 40238 43374 40290 43426
rect 47294 43374 47346 43426
rect 6974 43262 7026 43314
rect 7758 43262 7810 43314
rect 23550 43262 23602 43314
rect 34190 43262 34242 43314
rect 35422 43262 35474 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 28702 42926 28754 42978
rect 29934 42926 29986 42978
rect 30382 42926 30434 42978
rect 34526 42926 34578 42978
rect 2830 42814 2882 42866
rect 3278 42814 3330 42866
rect 7310 42814 7362 42866
rect 9998 42814 10050 42866
rect 15262 42814 15314 42866
rect 17390 42814 17442 42866
rect 20862 42814 20914 42866
rect 21646 42814 21698 42866
rect 23774 42814 23826 42866
rect 25118 42814 25170 42866
rect 27246 42814 27298 42866
rect 30158 42814 30210 42866
rect 30606 42814 30658 42866
rect 34414 42814 34466 42866
rect 4174 42702 4226 42754
rect 12910 42702 12962 42754
rect 13694 42702 13746 42754
rect 14030 42702 14082 42754
rect 14478 42702 14530 42754
rect 17950 42702 18002 42754
rect 24558 42702 24610 42754
rect 27918 42702 27970 42754
rect 28590 42702 28642 42754
rect 32846 42702 32898 42754
rect 8206 42590 8258 42642
rect 9102 42590 9154 42642
rect 12126 42590 12178 42642
rect 18734 42590 18786 42642
rect 31390 42590 31442 42642
rect 31502 42590 31554 42642
rect 31614 42590 31666 42642
rect 33070 42590 33122 42642
rect 33742 42590 33794 42642
rect 33966 42590 34018 42642
rect 1822 42478 1874 42530
rect 3726 42478 3778 42530
rect 4622 42478 4674 42530
rect 5070 42478 5122 42530
rect 5854 42478 5906 42530
rect 6302 42478 6354 42530
rect 6750 42478 6802 42530
rect 7758 42478 7810 42530
rect 8542 42478 8594 42530
rect 9214 42478 9266 42530
rect 9326 42478 9378 42530
rect 13806 42478 13858 42530
rect 28702 42478 28754 42530
rect 29486 42478 29538 42530
rect 31166 42478 31218 42530
rect 31278 42478 31330 42530
rect 32510 42478 32562 42530
rect 33854 42478 33906 42530
rect 34862 42478 34914 42530
rect 35310 42478 35362 42530
rect 36206 42814 36258 42866
rect 37998 42814 38050 42866
rect 35758 42702 35810 42754
rect 36654 42702 36706 42754
rect 40126 42590 40178 42642
rect 35646 42478 35698 42530
rect 37438 42478 37490 42530
rect 38446 42478 38498 42530
rect 38782 42478 38834 42530
rect 39230 42478 39282 42530
rect 39678 42478 39730 42530
rect 40574 42478 40626 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 18286 42142 18338 42194
rect 34974 42142 35026 42194
rect 36878 42142 36930 42194
rect 38222 42142 38274 42194
rect 6974 42030 7026 42082
rect 7534 42030 7586 42082
rect 7870 42030 7922 42082
rect 8430 42030 8482 42082
rect 8990 42030 9042 42082
rect 9886 42030 9938 42082
rect 9998 42030 10050 42082
rect 22766 42030 22818 42082
rect 31950 42030 32002 42082
rect 34862 42030 34914 42082
rect 2158 41918 2210 41970
rect 5182 41918 5234 41970
rect 5742 41918 5794 41970
rect 6638 41918 6690 41970
rect 8654 41918 8706 41970
rect 10558 41918 10610 41970
rect 14142 41918 14194 41970
rect 14814 41918 14866 41970
rect 17838 41918 17890 41970
rect 18398 41918 18450 41970
rect 22094 41918 22146 41970
rect 24110 41918 24162 41970
rect 24334 41918 24386 41970
rect 25790 41918 25842 41970
rect 29822 41918 29874 41970
rect 30046 41918 30098 41970
rect 30382 41918 30434 41970
rect 30718 41918 30770 41970
rect 34190 41918 34242 41970
rect 37326 41918 37378 41970
rect 37774 41918 37826 41970
rect 2606 41806 2658 41858
rect 3054 41806 3106 41858
rect 3502 41806 3554 41858
rect 3950 41806 4002 41858
rect 4398 41806 4450 41858
rect 4846 41806 4898 41858
rect 6078 41806 6130 41858
rect 8878 41806 8930 41858
rect 11342 41806 11394 41858
rect 13470 41806 13522 41858
rect 16942 41806 16994 41858
rect 19182 41806 19234 41858
rect 21422 41806 21474 41858
rect 23214 41806 23266 41858
rect 26462 41806 26514 41858
rect 28590 41806 28642 41858
rect 30494 41806 30546 41858
rect 35534 41806 35586 41858
rect 35982 41806 36034 41858
rect 36430 41806 36482 41858
rect 38670 41806 38722 41858
rect 39118 41806 39170 41858
rect 39566 41806 39618 41858
rect 40014 41806 40066 41858
rect 40462 41806 40514 41858
rect 41470 41806 41522 41858
rect 5518 41694 5570 41746
rect 5854 41694 5906 41746
rect 6078 41694 6130 41746
rect 6302 41694 6354 41746
rect 9886 41694 9938 41746
rect 17950 41694 18002 41746
rect 18174 41694 18226 41746
rect 24446 41694 24498 41746
rect 29934 41694 29986 41746
rect 32062 41694 32114 41746
rect 32286 41694 32338 41746
rect 32510 41694 32562 41746
rect 32622 41694 32674 41746
rect 33630 41694 33682 41746
rect 33966 41694 34018 41746
rect 35086 41694 35138 41746
rect 35982 41694 36034 41746
rect 36766 41694 36818 41746
rect 38894 41694 38946 41746
rect 39678 41694 39730 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 2606 41358 2658 41410
rect 3054 41358 3106 41410
rect 2830 41246 2882 41298
rect 3278 41246 3330 41298
rect 4062 41246 4114 41298
rect 4510 41246 4562 41298
rect 9326 41246 9378 41298
rect 9998 41246 10050 41298
rect 14478 41246 14530 41298
rect 23662 41246 23714 41298
rect 25342 41246 25394 41298
rect 26910 41246 26962 41298
rect 29598 41246 29650 41298
rect 34414 41246 34466 41298
rect 34974 41246 35026 41298
rect 38782 41246 38834 41298
rect 39678 41246 39730 41298
rect 40574 41246 40626 41298
rect 2382 41134 2434 41186
rect 6078 41134 6130 41186
rect 7758 41134 7810 41186
rect 8654 41134 8706 41186
rect 8990 41134 9042 41186
rect 9438 41134 9490 41186
rect 12910 41134 12962 41186
rect 14590 41134 14642 41186
rect 15262 41134 15314 41186
rect 15598 41134 15650 41186
rect 17054 41134 17106 41186
rect 17502 41134 17554 41186
rect 18510 41134 18562 41186
rect 18958 41134 19010 41186
rect 19966 41134 20018 41186
rect 21758 41134 21810 41186
rect 22654 41134 22706 41186
rect 24222 41134 24274 41186
rect 24670 41134 24722 41186
rect 26686 41134 26738 41186
rect 27694 41134 27746 41186
rect 28254 41134 28306 41186
rect 31726 41134 31778 41186
rect 32398 41134 32450 41186
rect 33070 41134 33122 41186
rect 34638 41134 34690 41186
rect 36654 41134 36706 41186
rect 6638 41022 6690 41074
rect 6974 41022 7026 41074
rect 7534 41022 7586 41074
rect 12126 41022 12178 41074
rect 14030 41022 14082 41074
rect 16046 41022 16098 41074
rect 16718 41022 16770 41074
rect 20862 41022 20914 41074
rect 27022 41022 27074 41074
rect 33294 41022 33346 41074
rect 33406 41022 33458 41074
rect 33518 41022 33570 41074
rect 35870 41022 35922 41074
rect 38334 41022 38386 41074
rect 40126 41022 40178 41074
rect 1934 40910 1986 40962
rect 3726 40910 3778 40962
rect 5070 40910 5122 40962
rect 5742 40910 5794 40962
rect 8094 40910 8146 40962
rect 9214 40910 9266 40962
rect 13806 40910 13858 40962
rect 17838 40910 17890 40962
rect 20750 40910 20802 40962
rect 28702 40910 28754 40962
rect 33182 40910 33234 40962
rect 35534 40910 35586 40962
rect 36430 40910 36482 40962
rect 37438 40910 37490 40962
rect 37886 40910 37938 40962
rect 39230 40910 39282 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 2158 40574 2210 40626
rect 3502 40574 3554 40626
rect 5630 40574 5682 40626
rect 6078 40574 6130 40626
rect 9662 40574 9714 40626
rect 3054 40462 3106 40514
rect 6638 40462 6690 40514
rect 7534 40462 7586 40514
rect 8430 40462 8482 40514
rect 9886 40462 9938 40514
rect 9998 40518 10050 40570
rect 18174 40574 18226 40626
rect 19630 40574 19682 40626
rect 23550 40574 23602 40626
rect 31502 40574 31554 40626
rect 34750 40574 34802 40626
rect 35534 40574 35586 40626
rect 35982 40574 36034 40626
rect 37774 40574 37826 40626
rect 38222 40574 38274 40626
rect 22990 40462 23042 40514
rect 24446 40462 24498 40514
rect 26462 40462 26514 40514
rect 29262 40462 29314 40514
rect 30270 40462 30322 40514
rect 48078 40462 48130 40514
rect 3950 40350 4002 40402
rect 4398 40350 4450 40402
rect 6974 40350 7026 40402
rect 7870 40350 7922 40402
rect 10558 40350 10610 40402
rect 11342 40350 11394 40402
rect 14142 40350 14194 40402
rect 14814 40350 14866 40402
rect 17614 40350 17666 40402
rect 18062 40350 18114 40402
rect 18286 40350 18338 40402
rect 19182 40350 19234 40402
rect 19966 40350 20018 40402
rect 20750 40350 20802 40402
rect 21198 40350 21250 40402
rect 22206 40350 22258 40402
rect 22878 40350 22930 40402
rect 24558 40350 24610 40402
rect 25790 40350 25842 40402
rect 29374 40350 29426 40402
rect 30046 40350 30098 40402
rect 30942 40350 30994 40402
rect 32622 40350 32674 40402
rect 33966 40350 34018 40402
rect 34190 40350 34242 40402
rect 35086 40350 35138 40402
rect 36430 40350 36482 40402
rect 39118 40350 39170 40402
rect 39566 40350 39618 40402
rect 2606 40238 2658 40290
rect 4734 40238 4786 40290
rect 5294 40238 5346 40290
rect 13470 40238 13522 40290
rect 16942 40238 16994 40290
rect 18846 40238 18898 40290
rect 28590 40238 28642 40290
rect 32286 40238 32338 40290
rect 36878 40238 36930 40290
rect 37326 40238 37378 40290
rect 38670 40238 38722 40290
rect 3838 40126 3890 40178
rect 4734 40126 4786 40178
rect 5070 40126 5122 40178
rect 8654 40126 8706 40178
rect 8990 40126 9042 40178
rect 31950 40126 32002 40178
rect 32062 40126 32114 40178
rect 32510 40126 32562 40178
rect 33630 40126 33682 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 7086 39790 7138 39842
rect 7646 39790 7698 39842
rect 9102 39790 9154 39842
rect 28702 39790 28754 39842
rect 29598 39790 29650 39842
rect 29822 39790 29874 39842
rect 32510 39790 32562 39842
rect 34862 39790 34914 39842
rect 35198 39790 35250 39842
rect 1822 39678 1874 39730
rect 2382 39678 2434 39730
rect 2830 39678 2882 39730
rect 3614 39678 3666 39730
rect 4510 39678 4562 39730
rect 5630 39678 5682 39730
rect 6190 39678 6242 39730
rect 7086 39678 7138 39730
rect 8094 39678 8146 39730
rect 12910 39678 12962 39730
rect 14478 39678 14530 39730
rect 20862 39678 20914 39730
rect 24558 39678 24610 39730
rect 25118 39678 25170 39730
rect 31166 39678 31218 39730
rect 31390 39678 31442 39730
rect 33070 39678 33122 39730
rect 33742 39678 33794 39730
rect 35534 39678 35586 39730
rect 37886 39678 37938 39730
rect 3278 39566 3330 39618
rect 10110 39566 10162 39618
rect 17278 39566 17330 39618
rect 17950 39566 18002 39618
rect 21646 39566 21698 39618
rect 27918 39566 27970 39618
rect 28590 39566 28642 39618
rect 30158 39566 30210 39618
rect 30270 39566 30322 39618
rect 31726 39566 31778 39618
rect 32846 39566 32898 39618
rect 33630 39566 33682 39618
rect 38334 39566 38386 39618
rect 38782 39566 38834 39618
rect 7982 39454 8034 39506
rect 8878 39454 8930 39506
rect 10782 39454 10834 39506
rect 13582 39454 13634 39506
rect 13918 39454 13970 39506
rect 16606 39454 16658 39506
rect 18734 39454 18786 39506
rect 22430 39454 22482 39506
rect 27246 39454 27298 39506
rect 33966 39454 34018 39506
rect 34638 39454 34690 39506
rect 35086 39454 35138 39506
rect 4174 39342 4226 39394
rect 5070 39342 5122 39394
rect 6526 39342 6578 39394
rect 7422 39342 7474 39394
rect 8206 39342 8258 39394
rect 9438 39342 9490 39394
rect 13806 39342 13858 39394
rect 28702 39342 28754 39394
rect 30382 39342 30434 39394
rect 30494 39342 30546 39394
rect 34526 39342 34578 39394
rect 35982 39342 36034 39394
rect 36430 39342 36482 39394
rect 37438 39342 37490 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 3726 39006 3778 39058
rect 5070 39006 5122 39058
rect 5854 39006 5906 39058
rect 7758 39006 7810 39058
rect 9102 39006 9154 39058
rect 10222 39006 10274 39058
rect 11790 39006 11842 39058
rect 33518 39006 33570 39058
rect 34414 39006 34466 39058
rect 35758 39006 35810 39058
rect 36206 39006 36258 39058
rect 36654 39006 36706 39058
rect 37102 39006 37154 39058
rect 1822 38894 1874 38946
rect 6414 38894 6466 38946
rect 14814 38894 14866 38946
rect 20414 38894 20466 38946
rect 21422 38894 21474 38946
rect 27806 38894 27858 38946
rect 29262 38894 29314 38946
rect 29486 38894 29538 38946
rect 29710 38894 29762 38946
rect 31278 38894 31330 38946
rect 32174 38894 32226 38946
rect 32846 38894 32898 38946
rect 37550 38894 37602 38946
rect 4174 38782 4226 38834
rect 10222 38782 10274 38834
rect 10334 38782 10386 38834
rect 10558 38782 10610 38834
rect 12910 38782 12962 38834
rect 14142 38782 14194 38834
rect 18286 38782 18338 38834
rect 19182 38782 19234 38834
rect 19742 38782 19794 38834
rect 20526 38782 20578 38834
rect 21086 38782 21138 38834
rect 21982 38782 22034 38834
rect 28478 38782 28530 38834
rect 30046 38782 30098 38834
rect 30158 38782 30210 38834
rect 31726 38782 31778 38834
rect 32398 38782 32450 38834
rect 33966 38782 34018 38834
rect 35310 38782 35362 38834
rect 4622 38670 4674 38722
rect 5518 38670 5570 38722
rect 6750 38670 6802 38722
rect 7310 38670 7362 38722
rect 8094 38670 8146 38722
rect 8542 38670 8594 38722
rect 11230 38670 11282 38722
rect 11454 38670 11506 38722
rect 13022 38670 13074 38722
rect 13358 38670 13410 38722
rect 16942 38670 16994 38722
rect 17614 38670 17666 38722
rect 22766 38670 22818 38722
rect 24894 38670 24946 38722
rect 25678 38670 25730 38722
rect 29150 38670 29202 38722
rect 31950 38670 32002 38722
rect 34862 38670 34914 38722
rect 17614 38558 17666 38610
rect 17950 38558 18002 38610
rect 30718 38558 30770 38610
rect 31054 38558 31106 38610
rect 32510 38558 32562 38610
rect 32734 38558 32786 38610
rect 33518 38558 33570 38610
rect 34190 38558 34242 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 6862 38222 6914 38274
rect 7534 38222 7586 38274
rect 7758 38222 7810 38274
rect 8206 38222 8258 38274
rect 12350 38222 12402 38274
rect 30158 38222 30210 38274
rect 32174 38222 32226 38274
rect 32398 38222 32450 38274
rect 33182 38222 33234 38274
rect 34078 38222 34130 38274
rect 35758 38222 35810 38274
rect 36654 38222 36706 38274
rect 4062 38110 4114 38162
rect 4622 38110 4674 38162
rect 5854 38110 5906 38162
rect 6638 38110 6690 38162
rect 9886 38110 9938 38162
rect 17390 38110 17442 38162
rect 20862 38110 20914 38162
rect 24558 38110 24610 38162
rect 28030 38110 28082 38162
rect 33070 38110 33122 38162
rect 36206 38110 36258 38162
rect 10670 37998 10722 38050
rect 12126 37998 12178 38050
rect 12574 37998 12626 38050
rect 12798 37998 12850 38050
rect 14030 37998 14082 38050
rect 14590 37998 14642 38050
rect 17950 37998 18002 38050
rect 21646 37998 21698 38050
rect 25230 37998 25282 38050
rect 29822 37998 29874 38050
rect 30942 37998 30994 38050
rect 32622 37998 32674 38050
rect 35758 37998 35810 38050
rect 5070 37886 5122 37938
rect 7534 37886 7586 37938
rect 7982 37886 8034 37938
rect 8430 37886 8482 37938
rect 10334 37886 10386 37938
rect 13694 37886 13746 37938
rect 15262 37886 15314 37938
rect 18734 37886 18786 37938
rect 22430 37886 22482 37938
rect 25902 37886 25954 37938
rect 28590 37886 28642 37938
rect 29598 37886 29650 37938
rect 30718 37886 30770 37938
rect 31278 37886 31330 37938
rect 31950 37886 32002 37938
rect 33966 37886 34018 37938
rect 6302 37774 6354 37826
rect 7198 37774 7250 37826
rect 8990 37774 9042 37826
rect 9326 37774 9378 37826
rect 11230 37774 11282 37826
rect 11566 37774 11618 37826
rect 12238 37774 12290 37826
rect 13806 37774 13858 37826
rect 28702 37774 28754 37826
rect 28926 37774 28978 37826
rect 30830 37774 30882 37826
rect 32062 37774 32114 37826
rect 33518 37774 33570 37826
rect 34414 37774 34466 37826
rect 34862 37774 34914 37826
rect 35310 37774 35362 37826
rect 36654 37774 36706 37826
rect 48078 37774 48130 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 5966 37438 6018 37490
rect 6302 37438 6354 37490
rect 7758 37438 7810 37490
rect 8654 37438 8706 37490
rect 9998 37438 10050 37490
rect 11454 37438 11506 37490
rect 12238 37438 12290 37490
rect 18062 37438 18114 37490
rect 31278 37438 31330 37490
rect 32734 37438 32786 37490
rect 34862 37438 34914 37490
rect 1822 37326 1874 37378
rect 16158 37326 16210 37378
rect 18398 37326 18450 37378
rect 18622 37326 18674 37378
rect 23886 37326 23938 37378
rect 25902 37326 25954 37378
rect 27246 37326 27298 37378
rect 28702 37326 28754 37378
rect 29262 37326 29314 37378
rect 30158 37326 30210 37378
rect 30382 37326 30434 37378
rect 33966 37326 34018 37378
rect 6862 37214 6914 37266
rect 11118 37214 11170 37266
rect 13470 37214 13522 37266
rect 16830 37214 16882 37266
rect 18958 37214 19010 37266
rect 22318 37214 22370 37266
rect 27022 37214 27074 37266
rect 28590 37214 28642 37266
rect 28814 37214 28866 37266
rect 29710 37214 29762 37266
rect 30942 37214 30994 37266
rect 33518 37214 33570 37266
rect 5518 37102 5570 37154
rect 7198 37102 7250 37154
rect 8206 37102 8258 37154
rect 8990 37102 9042 37154
rect 10446 37102 10498 37154
rect 12350 37102 12402 37154
rect 14030 37102 14082 37154
rect 19518 37102 19570 37154
rect 21646 37102 21698 37154
rect 23998 37102 24050 37154
rect 25678 37102 25730 37154
rect 29934 37102 29986 37154
rect 31726 37102 31778 37154
rect 32174 37102 32226 37154
rect 34414 37102 34466 37154
rect 35310 37102 35362 37154
rect 35758 37102 35810 37154
rect 10558 36990 10610 37042
rect 12014 36990 12066 37042
rect 12910 36990 12962 37042
rect 13246 36990 13298 37042
rect 23102 36990 23154 37042
rect 35310 36990 35362 37042
rect 35646 36990 35698 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 6974 36654 7026 36706
rect 7646 36654 7698 36706
rect 8990 36654 9042 36706
rect 9326 36654 9378 36706
rect 26126 36654 26178 36706
rect 30382 36654 30434 36706
rect 31390 36654 31442 36706
rect 34638 36654 34690 36706
rect 34862 36654 34914 36706
rect 6302 36542 6354 36594
rect 7646 36542 7698 36594
rect 8430 36542 8482 36594
rect 8878 36542 8930 36594
rect 10222 36542 10274 36594
rect 10670 36542 10722 36594
rect 15262 36542 15314 36594
rect 17390 36542 17442 36594
rect 17950 36542 18002 36594
rect 21646 36542 21698 36594
rect 23774 36542 23826 36594
rect 26014 36542 26066 36594
rect 27470 36542 27522 36594
rect 31390 36542 31442 36594
rect 32734 36542 32786 36594
rect 34078 36542 34130 36594
rect 34862 36542 34914 36594
rect 14030 36430 14082 36482
rect 14590 36430 14642 36482
rect 20078 36430 20130 36482
rect 20750 36430 20802 36482
rect 24446 36430 24498 36482
rect 25342 36430 25394 36482
rect 27134 36430 27186 36482
rect 27246 36430 27298 36482
rect 28590 36430 28642 36482
rect 29598 36430 29650 36482
rect 30382 36430 30434 36482
rect 9326 36318 9378 36370
rect 11230 36318 11282 36370
rect 11678 36318 11730 36370
rect 12910 36318 12962 36370
rect 13694 36318 13746 36370
rect 13806 36318 13858 36370
rect 26798 36318 26850 36370
rect 27694 36318 27746 36370
rect 28254 36318 28306 36370
rect 28814 36318 28866 36370
rect 29934 36318 29986 36370
rect 31726 36318 31778 36370
rect 6750 36206 6802 36258
rect 7086 36206 7138 36258
rect 7982 36206 8034 36258
rect 9774 36206 9826 36258
rect 12014 36206 12066 36258
rect 12574 36206 12626 36258
rect 27806 36206 27858 36258
rect 28366 36206 28418 36258
rect 29822 36206 29874 36258
rect 30830 36206 30882 36258
rect 32174 36206 32226 36258
rect 33070 36206 33122 36258
rect 33630 36206 33682 36258
rect 34414 36206 34466 36258
rect 48078 36206 48130 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 8094 35870 8146 35922
rect 8990 35870 9042 35922
rect 10782 35870 10834 35922
rect 13582 35870 13634 35922
rect 14478 35870 14530 35922
rect 15486 35870 15538 35922
rect 16606 35870 16658 35922
rect 18846 35870 18898 35922
rect 22878 35870 22930 35922
rect 26462 35870 26514 35922
rect 27134 35870 27186 35922
rect 29150 35870 29202 35922
rect 30606 35870 30658 35922
rect 31950 35870 32002 35922
rect 32846 35870 32898 35922
rect 33518 35870 33570 35922
rect 1822 35758 1874 35810
rect 12574 35758 12626 35810
rect 14142 35758 14194 35810
rect 17726 35758 17778 35810
rect 20078 35758 20130 35810
rect 24222 35758 24274 35810
rect 25902 35758 25954 35810
rect 28254 35758 28306 35810
rect 28590 35758 28642 35810
rect 29262 35758 29314 35810
rect 32398 35758 32450 35810
rect 8654 35646 8706 35698
rect 13246 35646 13298 35698
rect 15038 35646 15090 35698
rect 15374 35646 15426 35698
rect 15598 35646 15650 35698
rect 16158 35646 16210 35698
rect 16382 35646 16434 35698
rect 16942 35646 16994 35698
rect 18174 35646 18226 35698
rect 19294 35646 19346 35698
rect 22878 35646 22930 35698
rect 23326 35646 23378 35698
rect 23998 35646 24050 35698
rect 25678 35646 25730 35698
rect 26350 35646 26402 35698
rect 26574 35646 26626 35698
rect 31502 35646 31554 35698
rect 7310 35534 7362 35586
rect 7758 35534 7810 35586
rect 9886 35534 9938 35586
rect 10222 35534 10274 35586
rect 11230 35534 11282 35586
rect 11678 35534 11730 35586
rect 12014 35534 12066 35586
rect 22206 35534 22258 35586
rect 24782 35534 24834 35586
rect 24894 35534 24946 35586
rect 27470 35534 27522 35586
rect 27694 35534 27746 35586
rect 29710 35534 29762 35586
rect 30158 35534 30210 35586
rect 31166 35534 31218 35586
rect 12686 35422 12738 35474
rect 16606 35422 16658 35474
rect 17950 35422 18002 35474
rect 18398 35422 18450 35474
rect 26126 35422 26178 35474
rect 30382 35422 30434 35474
rect 31838 35422 31890 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 9326 35086 9378 35138
rect 9774 35086 9826 35138
rect 11678 35086 11730 35138
rect 12014 35086 12066 35138
rect 16494 35086 16546 35138
rect 25454 35086 25506 35138
rect 25678 35086 25730 35138
rect 27918 35086 27970 35138
rect 30158 35086 30210 35138
rect 32734 35086 32786 35138
rect 8878 34974 8930 35026
rect 9326 34974 9378 35026
rect 9774 34974 9826 35026
rect 10334 34974 10386 35026
rect 12014 34974 12066 35026
rect 14926 34974 14978 35026
rect 15710 34974 15762 35026
rect 17950 34974 18002 35026
rect 21646 34974 21698 35026
rect 29934 34974 29986 35026
rect 30942 34974 30994 35026
rect 31390 34974 31442 35026
rect 31726 34974 31778 35026
rect 11230 34862 11282 34914
rect 11566 34862 11618 34914
rect 15822 34862 15874 34914
rect 16942 34862 16994 34914
rect 17166 34862 17218 34914
rect 17390 34862 17442 34914
rect 20750 34862 20802 34914
rect 24446 34862 24498 34914
rect 25230 34862 25282 34914
rect 25790 34862 25842 34914
rect 26798 34862 26850 34914
rect 28590 34862 28642 34914
rect 30494 34862 30546 34914
rect 13806 34750 13858 34802
rect 14142 34750 14194 34802
rect 14702 34750 14754 34802
rect 15598 34750 15650 34802
rect 16046 34750 16098 34802
rect 20078 34750 20130 34802
rect 23774 34750 23826 34802
rect 27022 34750 27074 34802
rect 27694 34750 27746 34802
rect 10670 34638 10722 34690
rect 12574 34638 12626 34690
rect 13022 34638 13074 34690
rect 14926 34638 14978 34690
rect 25342 34638 25394 34690
rect 26462 34638 26514 34690
rect 27806 34638 27858 34690
rect 28478 34638 28530 34690
rect 29598 34638 29650 34690
rect 32174 34638 32226 34690
rect 32734 34638 32786 34690
rect 48078 34638 48130 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 9774 34302 9826 34354
rect 10222 34302 10274 34354
rect 11006 34302 11058 34354
rect 11566 34302 11618 34354
rect 12014 34302 12066 34354
rect 12462 34302 12514 34354
rect 12910 34302 12962 34354
rect 13694 34302 13746 34354
rect 15038 34302 15090 34354
rect 15934 34302 15986 34354
rect 24670 34302 24722 34354
rect 26574 34302 26626 34354
rect 27470 34302 27522 34354
rect 28030 34302 28082 34354
rect 28478 34302 28530 34354
rect 29822 34302 29874 34354
rect 30382 34302 30434 34354
rect 30718 34302 30770 34354
rect 31166 34302 31218 34354
rect 16494 34190 16546 34242
rect 25678 34190 25730 34242
rect 26014 34190 26066 34242
rect 26910 34190 26962 34242
rect 27582 34190 27634 34242
rect 13246 34078 13298 34130
rect 14702 34078 14754 34130
rect 15598 34078 15650 34130
rect 16718 34078 16770 34130
rect 17054 34078 17106 34130
rect 18062 34078 18114 34130
rect 18286 34078 18338 34130
rect 19182 34078 19234 34130
rect 23102 34078 23154 34130
rect 24222 34078 24274 34130
rect 24446 34078 24498 34130
rect 24894 34078 24946 34130
rect 27918 34078 27970 34130
rect 29374 34078 29426 34130
rect 10558 33966 10610 34018
rect 14142 33966 14194 34018
rect 16606 33966 16658 34018
rect 19854 33966 19906 34018
rect 21982 33966 22034 34018
rect 23438 33966 23490 34018
rect 24782 33966 24834 34018
rect 17726 33854 17778 33906
rect 17838 33854 17890 33906
rect 18398 33854 18450 33906
rect 23550 33854 23602 33906
rect 28926 33966 28978 34018
rect 28926 33854 28978 33906
rect 30158 33854 30210 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 3502 33518 3554 33570
rect 4174 33518 4226 33570
rect 13694 33518 13746 33570
rect 15038 33518 15090 33570
rect 19406 33518 19458 33570
rect 23774 33518 23826 33570
rect 24558 33518 24610 33570
rect 27694 33518 27746 33570
rect 27918 33518 27970 33570
rect 3838 33406 3890 33458
rect 11006 33406 11058 33458
rect 11678 33406 11730 33458
rect 12126 33406 12178 33458
rect 12574 33406 12626 33458
rect 14142 33406 14194 33458
rect 15486 33406 15538 33458
rect 15822 33406 15874 33458
rect 18622 33406 18674 33458
rect 20078 33406 20130 33458
rect 20862 33406 20914 33458
rect 21870 33406 21922 33458
rect 24782 33406 24834 33458
rect 26350 33406 26402 33458
rect 26910 33406 26962 33458
rect 27470 33406 27522 33458
rect 27918 33406 27970 33458
rect 28814 33406 28866 33458
rect 29486 33406 29538 33458
rect 4734 33294 4786 33346
rect 15038 33294 15090 33346
rect 17390 33294 17442 33346
rect 19742 33294 19794 33346
rect 21982 33294 22034 33346
rect 22654 33294 22706 33346
rect 23326 33294 23378 33346
rect 23550 33294 23602 33346
rect 23886 33294 23938 33346
rect 25678 33294 25730 33346
rect 4398 33182 4450 33234
rect 14590 33182 14642 33234
rect 23214 33182 23266 33234
rect 24782 33182 24834 33234
rect 25454 33182 25506 33234
rect 28366 33182 28418 33234
rect 1822 33070 1874 33122
rect 13022 33070 13074 33122
rect 13582 33070 13634 33122
rect 16382 33070 16434 33122
rect 16718 33070 16770 33122
rect 17614 33070 17666 33122
rect 18286 33070 18338 33122
rect 18510 33070 18562 33122
rect 18734 33070 18786 33122
rect 26462 33070 26514 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 12574 32734 12626 32786
rect 14926 32734 14978 32786
rect 16158 32734 16210 32786
rect 16830 32734 16882 32786
rect 17054 32734 17106 32786
rect 18846 32734 18898 32786
rect 22206 32734 22258 32786
rect 22318 32734 22370 32786
rect 25678 32734 25730 32786
rect 26014 32734 26066 32786
rect 27022 32734 27074 32786
rect 27470 32734 27522 32786
rect 27918 32734 27970 32786
rect 28366 32734 28418 32786
rect 13582 32622 13634 32674
rect 16718 32622 16770 32674
rect 19406 32622 19458 32674
rect 21086 32622 21138 32674
rect 22430 32622 22482 32674
rect 22542 32622 22594 32674
rect 23550 32622 23602 32674
rect 23998 32622 24050 32674
rect 24558 32622 24610 32674
rect 24894 32622 24946 32674
rect 48078 32622 48130 32674
rect 15374 32510 15426 32562
rect 19742 32510 19794 32562
rect 20190 32510 20242 32562
rect 20974 32510 21026 32562
rect 22990 32510 23042 32562
rect 23774 32510 23826 32562
rect 12238 32398 12290 32450
rect 13134 32398 13186 32450
rect 14030 32398 14082 32450
rect 14478 32398 14530 32450
rect 15710 32398 15762 32450
rect 17726 32398 17778 32450
rect 18286 32398 18338 32450
rect 23662 32398 23714 32450
rect 26574 32398 26626 32450
rect 18510 32286 18562 32338
rect 19518 32286 19570 32338
rect 19966 32286 20018 32338
rect 20750 32286 20802 32338
rect 21310 32286 21362 32338
rect 21534 32286 21586 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 14254 31838 14306 31890
rect 15598 31838 15650 31890
rect 21870 31838 21922 31890
rect 22878 31838 22930 31890
rect 24670 31838 24722 31890
rect 25230 31838 25282 31890
rect 25678 31838 25730 31890
rect 27022 31838 27074 31890
rect 16382 31726 16434 31778
rect 18510 31726 18562 31778
rect 19182 31726 19234 31778
rect 20190 31726 20242 31778
rect 20302 31726 20354 31778
rect 21646 31726 21698 31778
rect 22654 31726 22706 31778
rect 26574 31726 26626 31778
rect 16046 31614 16098 31666
rect 18286 31614 18338 31666
rect 20414 31614 20466 31666
rect 23214 31614 23266 31666
rect 24110 31614 24162 31666
rect 14702 31502 14754 31554
rect 15150 31502 15202 31554
rect 16942 31502 16994 31554
rect 17278 31502 17330 31554
rect 17838 31502 17890 31554
rect 19518 31502 19570 31554
rect 20862 31502 20914 31554
rect 22206 31502 22258 31554
rect 22990 31502 23042 31554
rect 23774 31502 23826 31554
rect 26126 31502 26178 31554
rect 48078 31502 48130 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 14814 31166 14866 31218
rect 16606 31166 16658 31218
rect 17054 31166 17106 31218
rect 18510 31166 18562 31218
rect 19742 31166 19794 31218
rect 23326 31166 23378 31218
rect 23550 31166 23602 31218
rect 19070 31054 19122 31106
rect 19518 31054 19570 31106
rect 22990 31054 23042 31106
rect 15598 30942 15650 30994
rect 18174 30942 18226 30994
rect 21870 30942 21922 30994
rect 22766 30942 22818 30994
rect 16158 30830 16210 30882
rect 17726 30830 17778 30882
rect 22094 30830 22146 30882
rect 16158 30718 16210 30770
rect 16494 30718 16546 30770
rect 16718 30718 16770 30770
rect 19854 30718 19906 30770
rect 20414 30718 20466 30770
rect 20526 30718 20578 30770
rect 20750 30718 20802 30770
rect 20862 30718 20914 30770
rect 24894 31166 24946 31218
rect 25678 31166 25730 31218
rect 23998 31054 24050 31106
rect 24446 30830 24498 30882
rect 26126 30830 26178 30882
rect 21534 30718 21586 30770
rect 23326 30718 23378 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 22206 30382 22258 30434
rect 22766 30382 22818 30434
rect 23438 30382 23490 30434
rect 17278 30270 17330 30322
rect 17838 30270 17890 30322
rect 19630 30270 19682 30322
rect 23438 30270 23490 30322
rect 24334 30270 24386 30322
rect 16158 30158 16210 30210
rect 18286 30158 18338 30210
rect 19182 30158 19234 30210
rect 20078 30158 20130 30210
rect 23886 30158 23938 30210
rect 25118 30158 25170 30210
rect 20862 30046 20914 30098
rect 21982 30046 22034 30098
rect 1822 29934 1874 29986
rect 18734 29934 18786 29986
rect 20526 29934 20578 29986
rect 21646 29934 21698 29986
rect 22430 29934 22482 29986
rect 22878 29934 22930 29986
rect 24782 29934 24834 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 19182 29598 19234 29650
rect 19742 29598 19794 29650
rect 20750 29598 20802 29650
rect 21198 29598 21250 29650
rect 21982 29598 22034 29650
rect 22542 29598 22594 29650
rect 22990 29598 23042 29650
rect 23438 29598 23490 29650
rect 23886 29598 23938 29650
rect 48078 29486 48130 29538
rect 20302 29262 20354 29314
rect 21646 29262 21698 29314
rect 20302 29150 20354 29202
rect 20638 29150 20690 29202
rect 21982 29150 22034 29202
rect 22542 29150 22594 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 21982 28702 22034 28754
rect 22542 28702 22594 28754
rect 22990 28702 23042 28754
rect 1822 28366 1874 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 1822 26798 1874 26850
rect 48078 26798 48130 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 1822 24782 1874 24834
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 48078 23662 48130 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 3502 23326 3554 23378
rect 3054 23102 3106 23154
rect 2046 22990 2098 23042
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 48078 22094 48130 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 1822 21646 1874 21698
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 1822 18958 1874 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 48078 18510 48130 18562
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 1822 17502 1874 17554
rect 48078 17390 48130 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 1822 15822 1874 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 1822 14254 1874 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 48078 12798 48130 12850
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 48078 12238 48130 12290
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 1822 10670 1874 10722
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 9102 9662 9154 9714
rect 8766 9550 8818 9602
rect 9550 9550 9602 9602
rect 48078 9550 48130 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 1822 9102 1874 9154
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 48078 7982 48130 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 1822 7534 1874 7586
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 48078 6414 48130 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 1822 4398 1874 4450
rect 2494 4398 2546 4450
rect 48078 4398 48130 4450
rect 47518 4174 47570 4226
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 4286 3614 4338 3666
rect 2158 3502 2210 3554
rect 3054 3502 3106 3554
rect 11902 3390 11954 3442
rect 12350 3390 12402 3442
rect 18622 3390 18674 3442
rect 19070 3390 19122 3442
rect 36430 3390 36482 3442
rect 37550 3390 37602 3442
rect 48078 3390 48130 3442
rect 3614 3278 3666 3330
rect 5742 3278 5794 3330
rect 9662 3278 9714 3330
rect 12686 3278 12738 3330
rect 14366 3278 14418 3330
rect 15710 3278 15762 3330
rect 17726 3278 17778 3330
rect 19406 3278 19458 3330
rect 21422 3278 21474 3330
rect 23102 3278 23154 3330
rect 26462 3278 26514 3330
rect 29262 3278 29314 3330
rect 31838 3278 31890 3330
rect 35198 3278 35250 3330
rect 37214 3278 37266 3330
rect 38558 3278 38610 3330
rect 41022 3278 41074 3330
rect 42590 3278 42642 3330
rect 43934 3278 43986 3330
rect 45950 3278 46002 3330
rect 47182 3278 47234 3330
rect 47742 3278 47794 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 40350 1822 40402 1874
rect 41022 1822 41074 1874
rect 8766 1710 8818 1762
rect 9662 1710 9714 1762
rect 20862 1710 20914 1762
rect 21422 1710 21474 1762
<< metal2 >>
rect 3276 49924 3332 49934
rect 672 49200 784 49800
rect 2016 49200 2128 49800
rect 700 47348 756 49200
rect 700 47282 756 47292
rect 1820 47796 1876 47806
rect 1820 45892 1876 47740
rect 2044 46450 2100 49200
rect 3164 49140 3220 49150
rect 2268 48356 2324 48366
rect 2044 46398 2046 46450
rect 2098 46398 2100 46450
rect 2044 46386 2100 46398
rect 2156 47124 2212 47134
rect 1820 45890 2100 45892
rect 1820 45838 1822 45890
rect 1874 45838 2100 45890
rect 1820 45836 2100 45838
rect 1820 45826 1876 45836
rect 1708 45780 1764 45790
rect 1708 45332 1764 45724
rect 1820 45332 1876 45342
rect 1708 45330 1876 45332
rect 1708 45278 1822 45330
rect 1874 45278 1876 45330
rect 1708 45276 1876 45278
rect 1820 45266 1876 45276
rect 1932 44996 1988 45006
rect 1932 43762 1988 44940
rect 1932 43710 1934 43762
rect 1986 43710 1988 43762
rect 1932 43698 1988 43710
rect 1820 42530 1876 42542
rect 1820 42478 1822 42530
rect 1874 42478 1876 42530
rect 1820 42420 1876 42478
rect 1820 42354 1876 42364
rect 2044 41524 2100 45836
rect 2156 45778 2212 47068
rect 2156 45726 2158 45778
rect 2210 45726 2212 45778
rect 2156 45714 2212 45726
rect 2156 44210 2212 44222
rect 2156 44158 2158 44210
rect 2210 44158 2212 44210
rect 2156 43764 2212 44158
rect 2156 43698 2212 43708
rect 2156 41972 2212 41982
rect 2156 41878 2212 41916
rect 1820 41468 2100 41524
rect 1820 39730 1876 41468
rect 2268 41188 2324 48300
rect 2492 47348 2548 47358
rect 2492 45330 2548 47292
rect 2716 46450 2772 46462
rect 2716 46398 2718 46450
rect 2770 46398 2772 46450
rect 2492 45278 2494 45330
rect 2546 45278 2548 45330
rect 2492 45266 2548 45278
rect 2604 45780 2660 45790
rect 2604 43708 2660 45724
rect 2716 45778 2772 46398
rect 2716 45726 2718 45778
rect 2770 45726 2772 45778
rect 2716 45714 2772 45726
rect 3164 45330 3220 49084
rect 3164 45278 3166 45330
rect 3218 45278 3220 45330
rect 3164 45266 3220 45278
rect 2492 43652 2660 43708
rect 3052 44322 3108 44334
rect 3052 44270 3054 44322
rect 3106 44270 3108 44322
rect 2380 43426 2436 43438
rect 2380 43374 2382 43426
rect 2434 43374 2436 43426
rect 2380 42084 2436 43374
rect 2380 42018 2436 42028
rect 2380 41188 2436 41198
rect 2268 41132 2380 41188
rect 2380 41094 2436 41132
rect 1820 39678 1822 39730
rect 1874 39678 1876 39730
rect 1820 39666 1876 39678
rect 1932 40964 1988 40974
rect 1820 38946 1876 38958
rect 1820 38894 1822 38946
rect 1874 38894 1876 38946
rect 1820 38388 1876 38894
rect 1820 38322 1876 38332
rect 1820 37378 1876 37390
rect 1820 37326 1822 37378
rect 1874 37326 1876 37378
rect 1820 37044 1876 37326
rect 1820 36978 1876 36988
rect 1820 35810 1876 35822
rect 1820 35758 1822 35810
rect 1874 35758 1876 35810
rect 1820 35028 1876 35758
rect 1820 34962 1876 34972
rect 1820 33122 1876 33134
rect 1820 33070 1822 33122
rect 1874 33070 1876 33122
rect 1820 33012 1876 33070
rect 1820 32946 1876 32956
rect 1820 29986 1876 29998
rect 1820 29934 1822 29986
rect 1874 29934 1876 29986
rect 1820 29652 1876 29934
rect 1820 29586 1876 29596
rect 1820 28418 1876 28430
rect 1820 28366 1822 28418
rect 1874 28366 1876 28418
rect 1820 28308 1876 28366
rect 1820 28242 1876 28252
rect 1820 26850 1876 26862
rect 1820 26798 1822 26850
rect 1874 26798 1876 26850
rect 1820 26292 1876 26798
rect 1820 26226 1876 26236
rect 1820 24834 1876 24846
rect 1820 24782 1822 24834
rect 1874 24782 1876 24834
rect 1820 24276 1876 24782
rect 1820 24210 1876 24220
rect 1932 23380 1988 40908
rect 2492 40740 2548 43652
rect 2716 43428 2772 43438
rect 2716 42196 2772 43372
rect 2828 43428 2884 43438
rect 3052 43428 3108 44270
rect 3164 43428 3220 43438
rect 2828 43426 2996 43428
rect 2828 43374 2830 43426
rect 2882 43374 2996 43426
rect 2828 43372 2996 43374
rect 2828 43362 2884 43372
rect 2828 42868 2884 42878
rect 2828 42774 2884 42812
rect 2716 42130 2772 42140
rect 2604 41860 2660 41870
rect 2604 41858 2772 41860
rect 2604 41806 2606 41858
rect 2658 41806 2772 41858
rect 2604 41804 2772 41806
rect 2604 41794 2660 41804
rect 2156 40684 2548 40740
rect 2604 41410 2660 41422
rect 2604 41358 2606 41410
rect 2658 41358 2660 41410
rect 2156 40626 2212 40684
rect 2156 40574 2158 40626
rect 2210 40574 2212 40626
rect 2156 40562 2212 40574
rect 2604 40516 2660 41358
rect 2492 40460 2660 40516
rect 2380 40404 2436 40414
rect 2380 39730 2436 40348
rect 2380 39678 2382 39730
rect 2434 39678 2436 39730
rect 2380 39666 2436 39678
rect 2492 39172 2548 40460
rect 2492 39106 2548 39116
rect 2604 40290 2660 40302
rect 2604 40238 2606 40290
rect 2658 40238 2660 40290
rect 2604 36148 2660 40238
rect 2716 37380 2772 41804
rect 2828 41748 2884 41758
rect 2828 41298 2884 41692
rect 2828 41246 2830 41298
rect 2882 41246 2884 41298
rect 2828 41234 2884 41246
rect 2828 39732 2884 39742
rect 2828 39638 2884 39676
rect 2940 38276 2996 43372
rect 3052 43426 3220 43428
rect 3052 43374 3166 43426
rect 3218 43374 3220 43426
rect 3052 43372 3220 43374
rect 3052 42644 3108 43372
rect 3164 43362 3220 43372
rect 3276 42866 3332 49868
rect 12236 49924 12292 49934
rect 4032 49200 4144 49800
rect 6048 49200 6160 49800
rect 6972 49252 7028 49262
rect 3836 48020 3892 48030
rect 3724 44884 3780 44894
rect 3724 44434 3780 44828
rect 3724 44382 3726 44434
rect 3778 44382 3780 44434
rect 3724 44370 3780 44382
rect 3724 43652 3780 43662
rect 3836 43652 3892 47964
rect 4060 46002 4116 49200
rect 7392 49200 7504 49800
rect 8092 49588 8148 49598
rect 5180 49028 5236 49038
rect 4956 48692 5012 48702
rect 4956 47124 5012 48636
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 4060 45950 4062 46002
rect 4114 45950 4116 46002
rect 4060 45938 4116 45950
rect 4844 45890 4900 45902
rect 4844 45838 4846 45890
rect 4898 45838 4900 45890
rect 4284 45332 4340 45342
rect 4172 44996 4228 45006
rect 3724 43650 3892 43652
rect 3724 43598 3726 43650
rect 3778 43598 3892 43650
rect 3724 43596 3892 43598
rect 4060 44994 4228 44996
rect 4060 44942 4174 44994
rect 4226 44942 4228 44994
rect 4060 44940 4228 44942
rect 3724 43586 3780 43596
rect 3276 42814 3278 42866
rect 3330 42814 3332 42866
rect 3276 42802 3332 42814
rect 3388 43316 3444 43326
rect 3052 42588 3332 42644
rect 3164 42196 3220 42206
rect 3052 41858 3108 41870
rect 3052 41806 3054 41858
rect 3106 41806 3108 41858
rect 3052 41410 3108 41806
rect 3052 41358 3054 41410
rect 3106 41358 3108 41410
rect 3052 41346 3108 41358
rect 3164 41300 3220 42140
rect 3276 41524 3332 42588
rect 3276 41458 3332 41468
rect 3276 41300 3332 41310
rect 3164 41298 3332 41300
rect 3164 41246 3278 41298
rect 3330 41246 3332 41298
rect 3164 41244 3332 41246
rect 3276 41234 3332 41244
rect 3388 41076 3444 43260
rect 4060 42980 4116 44940
rect 4172 44930 4228 44940
rect 4172 44436 4228 44446
rect 4284 44436 4340 45276
rect 4620 45332 4676 45342
rect 4620 45238 4676 45276
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4228 44380 4340 44436
rect 4172 44304 4228 44380
rect 4620 44324 4676 44334
rect 4620 44230 4676 44268
rect 4284 44212 4340 44222
rect 4172 43540 4228 43550
rect 4172 43446 4228 43484
rect 4060 42914 4116 42924
rect 4172 42756 4228 42766
rect 4172 42662 4228 42700
rect 3724 42532 3780 42542
rect 3724 42438 3780 42476
rect 3612 42084 3668 42094
rect 3500 41860 3556 41870
rect 3500 41766 3556 41804
rect 3276 41020 3444 41076
rect 3052 40516 3108 40526
rect 3052 40422 3108 40460
rect 3276 40068 3332 41020
rect 3612 40740 3668 42028
rect 3948 41858 4004 41870
rect 3948 41806 3950 41858
rect 4002 41806 4004 41858
rect 3948 41300 4004 41806
rect 3948 41234 4004 41244
rect 4060 41412 4116 41422
rect 4060 41298 4116 41356
rect 4060 41246 4062 41298
rect 4114 41246 4116 41298
rect 3724 40964 3780 40974
rect 3724 40962 3892 40964
rect 3724 40910 3726 40962
rect 3778 40910 3892 40962
rect 3724 40908 3892 40910
rect 3724 40898 3780 40908
rect 3612 40684 3780 40740
rect 3500 40628 3556 40638
rect 3500 40534 3556 40572
rect 2940 38210 2996 38220
rect 3164 40012 3332 40068
rect 3612 40292 3668 40302
rect 2716 37314 2772 37324
rect 2604 36082 2660 36092
rect 3164 31948 3220 40012
rect 3612 39732 3668 40236
rect 3276 39620 3332 39630
rect 3612 39600 3668 39676
rect 3276 39526 3332 39564
rect 3724 39058 3780 40684
rect 3836 40178 3892 40908
rect 3836 40126 3838 40178
rect 3890 40126 3892 40178
rect 3836 40114 3892 40126
rect 3948 40740 4004 40750
rect 3948 40402 4004 40684
rect 3948 40350 3950 40402
rect 4002 40350 4004 40402
rect 3724 39006 3726 39058
rect 3778 39006 3780 39058
rect 3724 38994 3780 39006
rect 3948 38836 4004 40350
rect 4060 40404 4116 41246
rect 4060 40338 4116 40348
rect 4284 41300 4340 44156
rect 4620 43426 4676 43438
rect 4620 43374 4622 43426
rect 4674 43374 4676 43426
rect 4620 43316 4676 43374
rect 4620 43250 4676 43260
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4620 42530 4676 42542
rect 4620 42478 4622 42530
rect 4674 42478 4676 42530
rect 4620 42420 4676 42478
rect 4620 42354 4676 42364
rect 4844 42084 4900 45838
rect 4956 44212 5012 47068
rect 5068 48132 5124 48142
rect 5068 45330 5124 48076
rect 5068 45278 5070 45330
rect 5122 45278 5124 45330
rect 5068 45266 5124 45278
rect 5068 44436 5124 44446
rect 5180 44436 5236 48972
rect 5964 48916 6020 48926
rect 5852 46452 5908 46462
rect 5852 46002 5908 46396
rect 5852 45950 5854 46002
rect 5906 45950 5908 46002
rect 5852 45938 5908 45950
rect 5964 45330 6020 48860
rect 6860 47796 6916 47806
rect 5964 45278 5966 45330
rect 6018 45278 6020 45330
rect 5516 44994 5572 45006
rect 5516 44942 5518 44994
rect 5570 44942 5572 44994
rect 5516 44660 5572 44942
rect 5516 44594 5572 44604
rect 5068 44434 5236 44436
rect 5068 44382 5070 44434
rect 5122 44382 5236 44434
rect 5068 44380 5236 44382
rect 5068 44370 5124 44380
rect 4956 44146 5012 44156
rect 4956 43652 5012 43662
rect 4956 43558 5012 43596
rect 5068 42530 5124 42542
rect 5068 42478 5070 42530
rect 5122 42478 5124 42530
rect 4844 42028 5012 42084
rect 4396 41860 4452 41870
rect 4396 41766 4452 41804
rect 4844 41858 4900 41870
rect 4844 41806 4846 41858
rect 4898 41806 4900 41858
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4508 41300 4564 41310
rect 4284 41298 4564 41300
rect 4284 41246 4510 41298
rect 4562 41246 4564 41298
rect 4284 41244 4564 41246
rect 4172 39394 4228 39406
rect 4172 39342 4174 39394
rect 4226 39342 4228 39394
rect 4172 39284 4228 39342
rect 4172 39218 4228 39228
rect 3724 38780 4004 38836
rect 4172 38836 4228 38846
rect 1932 23314 1988 23324
rect 2940 31892 3220 31948
rect 3500 33570 3556 33582
rect 3500 33518 3502 33570
rect 3554 33518 3556 33570
rect 2044 23042 2100 23054
rect 2044 22990 2046 23042
rect 2098 22990 2100 23042
rect 2044 22932 2100 22990
rect 2044 22866 2100 22876
rect 1820 21698 1876 21710
rect 1820 21646 1822 21698
rect 1874 21646 1876 21698
rect 1820 20916 1876 21646
rect 1820 20850 1876 20860
rect 2940 20132 2996 31892
rect 3500 23378 3556 33518
rect 3724 26908 3780 38780
rect 4172 38742 4228 38780
rect 4060 38164 4116 38174
rect 4060 38070 4116 38108
rect 4284 33908 4340 41244
rect 4508 41234 4564 41244
rect 4396 40404 4452 40414
rect 4396 40310 4452 40348
rect 4732 40290 4788 40302
rect 4732 40238 4734 40290
rect 4786 40238 4788 40290
rect 4732 40178 4788 40238
rect 4732 40126 4734 40178
rect 4786 40126 4788 40178
rect 4732 40114 4788 40126
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4508 39732 4564 39742
rect 4508 39638 4564 39676
rect 4620 38724 4676 38734
rect 4844 38724 4900 41806
rect 4620 38722 4900 38724
rect 4620 38670 4622 38722
rect 4674 38670 4900 38722
rect 4620 38668 4900 38670
rect 4620 38658 4676 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 4620 38276 4676 38286
rect 4620 38162 4676 38220
rect 4620 38110 4622 38162
rect 4674 38110 4676 38162
rect 4620 38098 4676 38110
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4844 36708 4900 38668
rect 4956 38164 5012 42028
rect 5068 41188 5124 42478
rect 5180 41970 5236 44380
rect 5852 44212 5908 44222
rect 5852 44118 5908 44156
rect 5964 43708 6020 45278
rect 5740 43652 6020 43708
rect 6076 47684 6132 47694
rect 6076 43708 6132 47628
rect 6524 47124 6580 47134
rect 6188 45668 6244 45678
rect 6188 45666 6356 45668
rect 6188 45614 6190 45666
rect 6242 45614 6356 45666
rect 6188 45612 6356 45614
rect 6188 45602 6244 45612
rect 6300 45108 6356 45612
rect 6300 44994 6356 45052
rect 6300 44942 6302 44994
rect 6354 44942 6356 44994
rect 6188 44100 6244 44110
rect 6300 44100 6356 44942
rect 6188 44098 6300 44100
rect 6188 44046 6190 44098
rect 6242 44046 6300 44098
rect 6188 44044 6300 44046
rect 6188 44034 6244 44044
rect 6076 43652 6244 43708
rect 5516 43426 5572 43438
rect 5516 43374 5518 43426
rect 5570 43374 5572 43426
rect 5516 43316 5572 43374
rect 5516 43250 5572 43260
rect 5180 41918 5182 41970
rect 5234 41918 5236 41970
rect 5180 41906 5236 41918
rect 5740 41970 5796 43652
rect 5964 43426 6020 43438
rect 5964 43374 5966 43426
rect 6018 43374 6020 43426
rect 5740 41918 5742 41970
rect 5794 41918 5796 41970
rect 5740 41906 5796 41918
rect 5852 42530 5908 42542
rect 5852 42478 5854 42530
rect 5906 42478 5908 42530
rect 5516 41746 5572 41758
rect 5516 41694 5518 41746
rect 5570 41694 5572 41746
rect 5068 41132 5460 41188
rect 5068 40962 5124 40974
rect 5068 40910 5070 40962
rect 5122 40910 5124 40962
rect 5068 40852 5124 40910
rect 5068 40786 5124 40796
rect 5292 40290 5348 40302
rect 5292 40238 5294 40290
rect 5346 40238 5348 40290
rect 5068 40178 5124 40190
rect 5068 40126 5070 40178
rect 5122 40126 5124 40178
rect 5068 39732 5124 40126
rect 5068 39666 5124 39676
rect 5068 39396 5124 39406
rect 5068 39394 5236 39396
rect 5068 39342 5070 39394
rect 5122 39342 5236 39394
rect 5068 39340 5236 39342
rect 5068 39330 5124 39340
rect 5068 39060 5124 39070
rect 5068 38966 5124 39004
rect 4956 38098 5012 38108
rect 5068 37940 5124 37950
rect 5068 37846 5124 37884
rect 4844 36642 4900 36652
rect 5180 36036 5236 39340
rect 5180 35970 5236 35980
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 5292 34580 5348 40238
rect 5404 39508 5460 41132
rect 5516 39956 5572 41694
rect 5852 41746 5908 42478
rect 5852 41694 5854 41746
rect 5906 41694 5908 41746
rect 5852 41682 5908 41694
rect 5964 41748 6020 43374
rect 6188 41972 6244 43652
rect 5964 41682 6020 41692
rect 6076 41858 6132 41870
rect 6076 41806 6078 41858
rect 6130 41806 6132 41858
rect 6076 41746 6132 41806
rect 6076 41694 6078 41746
rect 6130 41694 6132 41746
rect 6076 41682 6132 41694
rect 5852 41468 6132 41524
rect 5628 41412 5684 41422
rect 5628 40626 5684 41356
rect 5628 40574 5630 40626
rect 5682 40574 5684 40626
rect 5628 40562 5684 40574
rect 5740 40962 5796 40974
rect 5740 40910 5742 40962
rect 5794 40910 5796 40962
rect 5628 39956 5684 39966
rect 5516 39900 5628 39956
rect 5628 39730 5684 39900
rect 5628 39678 5630 39730
rect 5682 39678 5684 39730
rect 5628 39666 5684 39678
rect 5404 39452 5684 39508
rect 5404 39284 5460 39294
rect 5404 37156 5460 39228
rect 5516 38724 5572 38734
rect 5516 38630 5572 38668
rect 5516 37156 5572 37166
rect 5404 37154 5572 37156
rect 5404 37102 5518 37154
rect 5570 37102 5572 37154
rect 5404 37100 5572 37102
rect 5292 34514 5348 34524
rect 4284 33852 4900 33908
rect 4284 33796 4340 33852
rect 3836 33740 4340 33796
rect 4476 33740 4740 33750
rect 3836 33458 3892 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4172 33572 4228 33582
rect 4172 33570 4452 33572
rect 4172 33518 4174 33570
rect 4226 33518 4452 33570
rect 4172 33516 4452 33518
rect 4172 33506 4228 33516
rect 3836 33406 3838 33458
rect 3890 33406 3892 33458
rect 3836 33394 3892 33406
rect 4396 33234 4452 33516
rect 4732 33348 4788 33358
rect 4844 33348 4900 33852
rect 4732 33346 4900 33348
rect 4732 33294 4734 33346
rect 4786 33294 4900 33346
rect 4732 33292 4900 33294
rect 4732 33282 4788 33292
rect 4396 33182 4398 33234
rect 4450 33182 4452 33234
rect 4396 33170 4452 33182
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 5516 29540 5572 37100
rect 5628 36820 5684 39452
rect 5740 38836 5796 40910
rect 5852 39844 5908 41468
rect 5852 39396 5908 39788
rect 5852 39330 5908 39340
rect 5964 41300 6020 41310
rect 5852 39172 5908 39182
rect 5852 39058 5908 39116
rect 5852 39006 5854 39058
rect 5906 39006 5908 39058
rect 5852 38994 5908 39006
rect 5740 38770 5796 38780
rect 5964 38668 6020 41244
rect 6076 41186 6132 41468
rect 6076 41134 6078 41186
rect 6130 41134 6132 41186
rect 6076 41122 6132 41134
rect 6076 40628 6132 40638
rect 6188 40628 6244 41916
rect 6300 43652 6356 44044
rect 6300 43426 6356 43596
rect 6300 43374 6302 43426
rect 6354 43374 6356 43426
rect 6300 42530 6356 43374
rect 6524 42868 6580 47068
rect 6636 45668 6692 45678
rect 6636 45666 6804 45668
rect 6636 45614 6638 45666
rect 6690 45614 6804 45666
rect 6636 45612 6804 45614
rect 6636 45602 6692 45612
rect 6748 45108 6804 45612
rect 6748 45014 6804 45052
rect 6748 44436 6804 44446
rect 6748 44342 6804 44380
rect 6636 43652 6692 43662
rect 6636 43540 6692 43596
rect 6860 43652 6916 47740
rect 6860 43586 6916 43596
rect 6748 43540 6804 43550
rect 6636 43538 6804 43540
rect 6636 43486 6750 43538
rect 6802 43486 6804 43538
rect 6636 43484 6804 43486
rect 6748 43474 6804 43484
rect 6972 43314 7028 49196
rect 7084 47572 7140 47582
rect 7084 44436 7140 47516
rect 7196 46676 7252 46686
rect 7196 46002 7252 46620
rect 7196 45950 7198 46002
rect 7250 45950 7252 46002
rect 7196 45938 7252 45950
rect 7308 46004 7364 46014
rect 7308 45220 7364 45948
rect 7420 45780 7476 49200
rect 7644 45780 7700 45790
rect 7420 45778 7700 45780
rect 7420 45726 7646 45778
rect 7698 45726 7700 45778
rect 7420 45724 7700 45726
rect 7644 45714 7700 45724
rect 7868 45220 7924 45230
rect 7308 45164 7476 45220
rect 7308 44994 7364 45006
rect 7308 44942 7310 44994
rect 7362 44942 7364 44994
rect 7308 44548 7364 44942
rect 7308 44482 7364 44492
rect 7196 44436 7252 44446
rect 7084 44434 7252 44436
rect 7084 44382 7198 44434
rect 7250 44382 7252 44434
rect 7084 44380 7252 44382
rect 7196 44370 7252 44380
rect 6972 43262 6974 43314
rect 7026 43262 7028 43314
rect 6972 43250 7028 43262
rect 7308 43426 7364 43438
rect 7308 43374 7310 43426
rect 7362 43374 7364 43426
rect 7308 43204 7364 43374
rect 7308 43138 7364 43148
rect 7084 42980 7140 42990
rect 6580 42812 6692 42868
rect 6524 42802 6580 42812
rect 6300 42478 6302 42530
rect 6354 42478 6356 42530
rect 6300 41746 6356 42478
rect 6636 42196 6692 42812
rect 6748 42532 6804 42542
rect 6748 42530 6916 42532
rect 6748 42478 6750 42530
rect 6802 42478 6916 42530
rect 6748 42476 6916 42478
rect 6748 42466 6804 42476
rect 6636 42140 6804 42196
rect 6636 41972 6692 41982
rect 6636 41878 6692 41916
rect 6748 41748 6804 42140
rect 6300 41694 6302 41746
rect 6354 41694 6356 41746
rect 6300 41682 6356 41694
rect 6636 41692 6804 41748
rect 6860 41972 6916 42476
rect 6972 42084 7028 42094
rect 6972 41990 7028 42028
rect 6636 41074 6692 41692
rect 6636 41022 6638 41074
rect 6690 41022 6692 41074
rect 6636 41010 6692 41022
rect 6860 40740 6916 41916
rect 6972 41076 7028 41086
rect 6972 40982 7028 41020
rect 6860 40674 6916 40684
rect 6076 40626 6244 40628
rect 6076 40574 6078 40626
rect 6130 40574 6244 40626
rect 6076 40572 6244 40574
rect 6076 40562 6132 40572
rect 6636 40514 6692 40526
rect 6636 40462 6638 40514
rect 6690 40462 6692 40514
rect 6076 40180 6132 40190
rect 6076 39060 6132 40124
rect 6636 40180 6692 40462
rect 6972 40402 7028 40414
rect 6972 40350 6974 40402
rect 7026 40350 7028 40402
rect 6972 40292 7028 40350
rect 6972 40226 7028 40236
rect 6636 40114 6692 40124
rect 7084 40068 7140 42924
rect 7308 42868 7364 42878
rect 7420 42868 7476 45164
rect 7756 44994 7812 45006
rect 7756 44942 7758 44994
rect 7810 44942 7812 44994
rect 7644 44098 7700 44110
rect 7644 44046 7646 44098
rect 7698 44046 7700 44098
rect 7644 43876 7700 44046
rect 7644 43810 7700 43820
rect 7756 43708 7812 44942
rect 7308 42866 7476 42868
rect 7308 42814 7310 42866
rect 7362 42814 7476 42866
rect 7308 42812 7476 42814
rect 7532 43652 7812 43708
rect 7308 42802 7364 42812
rect 7532 42644 7588 43652
rect 7756 43426 7812 43438
rect 7756 43374 7758 43426
rect 7810 43374 7812 43426
rect 7756 43314 7812 43374
rect 7756 43262 7758 43314
rect 7810 43262 7812 43314
rect 7756 43250 7812 43262
rect 7308 42588 7588 42644
rect 6972 40012 7140 40068
rect 7196 40740 7252 40750
rect 6188 39956 6244 39966
rect 6188 39730 6244 39900
rect 6188 39678 6190 39730
rect 6242 39678 6244 39730
rect 6188 39666 6244 39678
rect 6860 39732 6916 39742
rect 6524 39396 6580 39406
rect 6860 39396 6916 39676
rect 6524 39394 6860 39396
rect 6524 39342 6526 39394
rect 6578 39342 6860 39394
rect 6524 39340 6860 39342
rect 6524 39330 6580 39340
rect 6076 38994 6132 39004
rect 6524 39172 6580 39182
rect 6412 38948 6468 38958
rect 6412 38854 6468 38892
rect 6524 38724 6580 39116
rect 5964 38612 6244 38668
rect 5852 38388 5908 38398
rect 5852 38162 5908 38332
rect 5852 38110 5854 38162
rect 5906 38110 5908 38162
rect 5852 38098 5908 38110
rect 5964 37492 6020 37502
rect 6188 37492 6244 38612
rect 6524 38164 6580 38668
rect 6748 38724 6804 38734
rect 6860 38724 6916 39340
rect 6748 38722 6916 38724
rect 6748 38670 6750 38722
rect 6802 38670 6916 38722
rect 6748 38668 6916 38670
rect 6636 38164 6692 38174
rect 6524 38162 6692 38164
rect 6524 38110 6638 38162
rect 6690 38110 6692 38162
rect 6524 38108 6692 38110
rect 6636 38098 6692 38108
rect 6748 38052 6804 38668
rect 6748 37986 6804 37996
rect 6860 38274 6916 38286
rect 6860 38222 6862 38274
rect 6914 38222 6916 38274
rect 6300 37826 6356 37838
rect 6300 37774 6302 37826
rect 6354 37774 6356 37826
rect 6300 37716 6356 37774
rect 6300 37660 6468 37716
rect 6300 37492 6356 37502
rect 6188 37490 6356 37492
rect 6188 37438 6302 37490
rect 6354 37438 6356 37490
rect 6188 37436 6356 37438
rect 5964 37398 6020 37436
rect 6300 37426 6356 37436
rect 5628 35364 5684 36764
rect 5628 35298 5684 35308
rect 6300 36596 6356 36606
rect 5516 29474 5572 29484
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 6300 27860 6356 36540
rect 6412 36484 6468 37660
rect 6860 37268 6916 38222
rect 6860 37174 6916 37212
rect 6972 36706 7028 40012
rect 7084 39842 7140 39854
rect 7084 39790 7086 39842
rect 7138 39790 7140 39842
rect 7084 39730 7140 39790
rect 7084 39678 7086 39730
rect 7138 39678 7140 39730
rect 7084 39666 7140 39678
rect 7196 39508 7252 40684
rect 7084 39452 7252 39508
rect 7084 38668 7140 39452
rect 7308 38948 7364 42588
rect 7756 42532 7812 42542
rect 7868 42532 7924 45164
rect 7644 42530 7924 42532
rect 7644 42478 7758 42530
rect 7810 42478 7924 42530
rect 7644 42476 7924 42478
rect 7980 45108 8036 45118
rect 7532 42084 7588 42094
rect 7420 42082 7588 42084
rect 7420 42030 7534 42082
rect 7586 42030 7588 42082
rect 7420 42028 7588 42030
rect 7420 40740 7476 42028
rect 7532 42018 7588 42028
rect 7532 41074 7588 41086
rect 7532 41022 7534 41074
rect 7586 41022 7588 41074
rect 7532 40964 7588 41022
rect 7532 40898 7588 40908
rect 7420 40674 7476 40684
rect 7532 40514 7588 40526
rect 7532 40462 7534 40514
rect 7586 40462 7588 40514
rect 7420 39396 7476 39406
rect 7420 39302 7476 39340
rect 7308 38892 7476 38948
rect 7308 38724 7364 38734
rect 7084 38612 7252 38668
rect 7308 38630 7364 38668
rect 7196 38276 7252 38612
rect 7420 38276 7476 38892
rect 7196 38220 7364 38276
rect 7308 37940 7364 38220
rect 7420 38210 7476 38220
rect 7532 38274 7588 40462
rect 7644 39842 7700 42476
rect 7756 42466 7812 42476
rect 7868 42196 7924 42206
rect 7868 42082 7924 42140
rect 7868 42030 7870 42082
rect 7922 42030 7924 42082
rect 7868 42018 7924 42030
rect 7756 41972 7812 41982
rect 7756 41412 7812 41916
rect 7756 41356 7924 41412
rect 7756 41186 7812 41198
rect 7756 41134 7758 41186
rect 7810 41134 7812 41186
rect 7756 40740 7812 41134
rect 7868 40964 7924 41356
rect 7868 40898 7924 40908
rect 7756 40674 7812 40684
rect 7868 40402 7924 40414
rect 7868 40350 7870 40402
rect 7922 40350 7924 40402
rect 7644 39790 7646 39842
rect 7698 39790 7700 39842
rect 7644 39778 7700 39790
rect 7756 40180 7812 40190
rect 7532 38222 7534 38274
rect 7586 38222 7588 38274
rect 7532 38210 7588 38222
rect 7644 39620 7700 39630
rect 7644 39396 7700 39564
rect 7756 39508 7812 40124
rect 7868 40068 7924 40350
rect 7868 40002 7924 40012
rect 7980 39732 8036 45052
rect 8092 44434 8148 49532
rect 9408 49200 9520 49800
rect 10668 49700 10724 49710
rect 9324 48356 9380 48366
rect 8540 48020 8596 48030
rect 8428 47964 8540 48020
rect 8428 47796 8484 47964
rect 8540 47954 8596 47964
rect 8428 47730 8484 47740
rect 8764 47796 8820 47806
rect 8540 47236 8596 47246
rect 8316 47124 8372 47134
rect 8316 47010 8372 47068
rect 8316 46958 8318 47010
rect 8370 46958 8372 47010
rect 8316 46946 8372 46958
rect 8540 47010 8596 47180
rect 8540 46958 8542 47010
rect 8594 46958 8596 47010
rect 8540 46946 8596 46958
rect 8428 46900 8484 46910
rect 8316 46788 8372 46798
rect 8204 45668 8260 45678
rect 8204 45574 8260 45612
rect 8204 45332 8260 45342
rect 8316 45332 8372 46732
rect 8204 45330 8372 45332
rect 8204 45278 8206 45330
rect 8258 45278 8372 45330
rect 8204 45276 8372 45278
rect 8204 45266 8260 45276
rect 8092 44382 8094 44434
rect 8146 44382 8148 44434
rect 8092 44370 8148 44382
rect 8428 44324 8484 46844
rect 8316 44268 8484 44324
rect 8540 45668 8596 45678
rect 8540 45330 8596 45612
rect 8540 45278 8542 45330
rect 8594 45278 8596 45330
rect 8316 43876 8372 44268
rect 8428 44100 8484 44110
rect 8540 44100 8596 45278
rect 8484 44044 8596 44100
rect 8428 43968 8484 44044
rect 8316 43820 8484 43876
rect 8204 43652 8260 43662
rect 8204 43558 8260 43596
rect 8204 42644 8260 42654
rect 8204 42550 8260 42588
rect 8428 42082 8484 43820
rect 8652 43428 8708 43438
rect 8652 43334 8708 43372
rect 8428 42030 8430 42082
rect 8482 42030 8484 42082
rect 8428 42018 8484 42030
rect 8540 42530 8596 42542
rect 8540 42478 8542 42530
rect 8594 42478 8596 42530
rect 8092 40964 8148 40974
rect 8092 40962 8372 40964
rect 8092 40910 8094 40962
rect 8146 40910 8372 40962
rect 8092 40908 8372 40910
rect 8092 40898 8148 40908
rect 8092 39732 8148 39742
rect 7980 39730 8148 39732
rect 7980 39678 8094 39730
rect 8146 39678 8148 39730
rect 7980 39676 8148 39678
rect 8092 39666 8148 39676
rect 7980 39508 8036 39518
rect 7756 39506 8036 39508
rect 7756 39454 7982 39506
rect 8034 39454 8036 39506
rect 7756 39452 8036 39454
rect 7196 37828 7252 37838
rect 7196 37734 7252 37772
rect 7196 37156 7252 37166
rect 7308 37156 7364 37884
rect 7532 37940 7588 37950
rect 7532 37846 7588 37884
rect 7644 37716 7700 39340
rect 7868 39284 7924 39294
rect 7756 39060 7812 39070
rect 7756 38966 7812 39004
rect 7756 38724 7812 38734
rect 7756 38274 7812 38668
rect 7756 38222 7758 38274
rect 7810 38222 7812 38274
rect 7756 38210 7812 38222
rect 7252 37100 7364 37156
rect 7532 37660 7700 37716
rect 7756 38052 7812 38062
rect 7196 37062 7252 37100
rect 6972 36654 6974 36706
rect 7026 36654 7028 36706
rect 6972 36642 7028 36654
rect 6412 36418 6468 36428
rect 6748 36260 6804 36270
rect 6748 36166 6804 36204
rect 7084 36258 7140 36270
rect 7084 36206 7086 36258
rect 7138 36206 7140 36258
rect 7084 35028 7140 36206
rect 7084 34962 7140 34972
rect 7308 35588 7364 35598
rect 6300 27794 6356 27804
rect 6636 33572 6692 33582
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 3724 26852 4004 26908
rect 3500 23326 3502 23378
rect 3554 23326 3556 23378
rect 3052 23156 3108 23166
rect 3500 23156 3556 23326
rect 3052 23154 3556 23156
rect 3052 23102 3054 23154
rect 3106 23102 3556 23154
rect 3052 23100 3556 23102
rect 3052 23090 3108 23100
rect 2940 20066 2996 20076
rect 1820 19010 1876 19022
rect 1820 18958 1822 19010
rect 1874 18958 1876 19010
rect 1820 18900 1876 18958
rect 1820 18834 1876 18844
rect 3948 18340 4004 26852
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 3948 18274 4004 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1820 17556 1876 17566
rect 1820 17462 1876 17500
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 1820 15874 1876 15886
rect 1820 15822 1822 15874
rect 1874 15822 1876 15874
rect 1820 15540 1876 15822
rect 1820 15474 1876 15484
rect 6636 15092 6692 33516
rect 7308 23268 7364 35532
rect 7532 30548 7588 37660
rect 7756 37490 7812 37996
rect 7756 37438 7758 37490
rect 7810 37438 7812 37490
rect 7756 37426 7812 37438
rect 7868 37492 7924 39228
rect 7980 38724 8036 39452
rect 8204 39396 8260 39406
rect 8204 39302 8260 39340
rect 7980 38658 8036 38668
rect 8092 38722 8148 38734
rect 8092 38670 8094 38722
rect 8146 38670 8148 38722
rect 7980 37940 8036 37950
rect 8092 37940 8148 38670
rect 7980 37938 8092 37940
rect 7980 37886 7982 37938
rect 8034 37886 8092 37938
rect 7980 37884 8092 37886
rect 7980 37874 8036 37884
rect 8092 37874 8148 37884
rect 8204 38274 8260 38286
rect 8204 38222 8206 38274
rect 8258 38222 8260 38274
rect 8204 37716 8260 38222
rect 7868 37426 7924 37436
rect 8092 37660 8260 37716
rect 7980 37156 8036 37166
rect 7644 36706 7700 36718
rect 7644 36654 7646 36706
rect 7698 36654 7700 36706
rect 7644 36594 7700 36654
rect 7644 36542 7646 36594
rect 7698 36542 7700 36594
rect 7644 36530 7700 36542
rect 7980 36258 8036 37100
rect 8092 36932 8148 37660
rect 8204 37156 8260 37166
rect 8204 37062 8260 37100
rect 8092 36876 8260 36932
rect 7980 36206 7982 36258
rect 8034 36206 8036 36258
rect 7532 30482 7588 30492
rect 7756 35588 7812 35598
rect 7756 24164 7812 35532
rect 7980 33572 8036 36206
rect 8092 36596 8148 36606
rect 8092 35922 8148 36540
rect 8092 35870 8094 35922
rect 8146 35870 8148 35922
rect 8092 35858 8148 35870
rect 8204 35028 8260 36876
rect 8204 34962 8260 34972
rect 8316 33684 8372 40908
rect 8428 40516 8484 40526
rect 8428 40422 8484 40460
rect 8540 38948 8596 42478
rect 8764 42532 8820 47740
rect 9100 47348 9156 47358
rect 8876 46450 8932 46462
rect 8876 46398 8878 46450
rect 8930 46398 8932 46450
rect 8876 45778 8932 46398
rect 8876 45726 8878 45778
rect 8930 45726 8932 45778
rect 8876 45714 8932 45726
rect 9100 45330 9156 47292
rect 9100 45278 9102 45330
rect 9154 45278 9156 45330
rect 9100 45266 9156 45278
rect 8988 44100 9044 44110
rect 8988 44006 9044 44044
rect 9100 43428 9156 43438
rect 8764 42466 8820 42476
rect 8876 43426 9156 43428
rect 8876 43374 9102 43426
rect 9154 43374 9156 43426
rect 8876 43372 9156 43374
rect 8876 42084 8932 43372
rect 9100 43362 9156 43372
rect 9100 42644 9156 42654
rect 9100 42550 9156 42588
rect 8764 42028 8932 42084
rect 8988 42532 9044 42542
rect 8988 42082 9044 42476
rect 8988 42030 8990 42082
rect 9042 42030 9044 42082
rect 8652 41970 8708 41982
rect 8652 41918 8654 41970
rect 8706 41918 8708 41970
rect 8652 41412 8708 41918
rect 8652 41346 8708 41356
rect 8764 41972 8820 42028
rect 8988 42018 9044 42030
rect 9212 42530 9268 42542
rect 9212 42478 9214 42530
rect 9266 42478 9268 42530
rect 9212 42084 9268 42478
rect 9324 42532 9380 48300
rect 9436 46450 9492 49200
rect 9436 46398 9438 46450
rect 9490 46398 9492 46450
rect 9436 46386 9492 46398
rect 10556 47684 10612 47694
rect 10556 47236 10612 47628
rect 10332 46340 10388 46350
rect 9772 46228 9828 46238
rect 9772 46002 9828 46172
rect 9772 45950 9774 46002
rect 9826 45950 9828 46002
rect 9772 45938 9828 45950
rect 10332 45778 10388 46284
rect 10332 45726 10334 45778
rect 10386 45726 10388 45778
rect 10332 45714 10388 45726
rect 9884 45108 9940 45118
rect 9772 44994 9828 45006
rect 9772 44942 9774 44994
rect 9826 44942 9828 44994
rect 9772 44772 9828 44942
rect 9772 44706 9828 44716
rect 9772 44548 9828 44558
rect 9772 44434 9828 44492
rect 9772 44382 9774 44434
rect 9826 44382 9828 44434
rect 9324 42438 9380 42476
rect 9436 44098 9492 44110
rect 9436 44046 9438 44098
rect 9490 44046 9492 44098
rect 9212 42018 9268 42028
rect 8652 41188 8708 41198
rect 8652 41094 8708 41132
rect 8764 40740 8820 41916
rect 8876 41860 8932 41870
rect 9436 41860 9492 44046
rect 8876 41766 8932 41804
rect 9100 41804 9492 41860
rect 9548 41860 9604 41870
rect 9100 41524 9156 41804
rect 8652 40684 8820 40740
rect 8876 41468 9156 41524
rect 9436 41636 9492 41646
rect 8652 40404 8708 40684
rect 8876 40516 8932 41468
rect 8988 41300 9044 41310
rect 8988 41186 9044 41244
rect 9324 41300 9380 41310
rect 9324 41206 9380 41244
rect 8988 41134 8990 41186
rect 9042 41134 9044 41186
rect 8988 40740 9044 41134
rect 9100 41188 9156 41198
rect 9100 40964 9156 41132
rect 9436 41186 9492 41580
rect 9436 41134 9438 41186
rect 9490 41134 9492 41186
rect 9436 41122 9492 41134
rect 9212 40964 9268 40974
rect 9100 40962 9268 40964
rect 9100 40910 9214 40962
rect 9266 40910 9268 40962
rect 9100 40908 9268 40910
rect 9212 40898 9268 40908
rect 9436 40852 9492 40862
rect 9436 40740 9492 40796
rect 8988 40684 9492 40740
rect 8876 40460 9380 40516
rect 8652 40348 8820 40404
rect 8652 40180 8708 40190
rect 8652 40086 8708 40124
rect 8764 39396 8820 40348
rect 8764 39330 8820 39340
rect 8876 40292 8932 40302
rect 8876 39506 8932 40236
rect 8876 39454 8878 39506
rect 8930 39454 8932 39506
rect 8540 38892 8820 38948
rect 8540 38722 8596 38734
rect 8540 38670 8542 38722
rect 8594 38670 8596 38722
rect 8540 38164 8596 38670
rect 8540 38098 8596 38108
rect 8428 37940 8484 37950
rect 8428 37846 8484 37884
rect 8652 37604 8708 37614
rect 8652 37490 8708 37548
rect 8652 37438 8654 37490
rect 8706 37438 8708 37490
rect 8652 37426 8708 37438
rect 8428 36596 8484 36606
rect 8428 36502 8484 36540
rect 8652 35700 8708 35710
rect 8652 35606 8708 35644
rect 8764 34356 8820 38892
rect 8876 36596 8932 39454
rect 8988 40178 9044 40190
rect 8988 40126 8990 40178
rect 9042 40126 9044 40178
rect 8988 38668 9044 40126
rect 9100 39844 9156 39854
rect 9100 39750 9156 39788
rect 9100 39396 9156 39406
rect 9100 39058 9156 39340
rect 9100 39006 9102 39058
rect 9154 39006 9156 39058
rect 9100 38994 9156 39006
rect 9212 39060 9268 39070
rect 8988 38612 9156 38668
rect 8988 37826 9044 37838
rect 8988 37774 8990 37826
rect 9042 37774 9044 37826
rect 8988 37380 9044 37774
rect 8988 37314 9044 37324
rect 8988 37154 9044 37166
rect 8988 37102 8990 37154
rect 9042 37102 9044 37154
rect 8988 36706 9044 37102
rect 8988 36654 8990 36706
rect 9042 36654 9044 36706
rect 8988 36642 9044 36654
rect 8876 36464 8932 36540
rect 8988 36260 9044 36270
rect 8988 35922 9044 36204
rect 8988 35870 8990 35922
rect 9042 35870 9044 35922
rect 8988 35858 9044 35870
rect 8876 35028 8932 35038
rect 8876 34934 8932 34972
rect 8764 34290 8820 34300
rect 8316 33618 8372 33628
rect 7980 33506 8036 33516
rect 9100 31332 9156 38612
rect 9100 31266 9156 31276
rect 9212 29764 9268 39004
rect 9324 38668 9380 40460
rect 9436 39396 9492 39406
rect 9436 39302 9492 39340
rect 9324 38612 9492 38668
rect 9324 37940 9380 37950
rect 9324 37826 9380 37884
rect 9324 37774 9326 37826
rect 9378 37774 9380 37826
rect 9324 36706 9380 37774
rect 9324 36654 9326 36706
rect 9378 36654 9380 36706
rect 9324 36372 9380 36654
rect 9324 36278 9380 36316
rect 9324 35138 9380 35150
rect 9324 35086 9326 35138
rect 9378 35086 9380 35138
rect 9324 35026 9380 35086
rect 9324 34974 9326 35026
rect 9378 34974 9380 35026
rect 9324 34962 9380 34974
rect 9436 34468 9492 38612
rect 9548 35252 9604 41804
rect 9772 41860 9828 44382
rect 9884 43650 9940 45052
rect 10220 44994 10276 45006
rect 10220 44942 10222 44994
rect 10274 44942 10276 44994
rect 10220 44548 10276 44942
rect 10220 44482 10276 44492
rect 10444 44322 10500 44334
rect 10444 44270 10446 44322
rect 10498 44270 10500 44322
rect 10444 43708 10500 44270
rect 10556 43988 10612 47180
rect 10668 45330 10724 49644
rect 11424 49200 11536 49800
rect 11676 49252 11732 49262
rect 10668 45278 10670 45330
rect 10722 45278 10724 45330
rect 10668 45266 10724 45278
rect 10780 48916 10836 48926
rect 10668 44212 10724 44222
rect 10780 44212 10836 48860
rect 11116 48468 11172 48478
rect 10892 45892 10948 45902
rect 10892 44996 10948 45836
rect 11004 45780 11060 45790
rect 11004 45686 11060 45724
rect 11116 45444 11172 48412
rect 11452 45892 11508 49200
rect 11676 46116 11732 49196
rect 11676 46050 11732 46060
rect 11788 48132 11844 48142
rect 11788 45892 11844 48076
rect 12124 47012 12180 47022
rect 11452 45826 11508 45836
rect 11676 45836 11844 45892
rect 11900 46002 11956 46014
rect 11900 45950 11902 46002
rect 11954 45950 11956 46002
rect 11564 45778 11620 45790
rect 11564 45726 11566 45778
rect 11618 45726 11620 45778
rect 10892 44930 10948 44940
rect 11004 45388 11172 45444
rect 11228 45556 11284 45566
rect 10668 44210 10836 44212
rect 10668 44158 10670 44210
rect 10722 44158 10836 44210
rect 10668 44156 10836 44158
rect 10668 44146 10724 44156
rect 11004 44100 11060 45388
rect 11116 45220 11172 45230
rect 11116 45126 11172 45164
rect 11228 44434 11284 45500
rect 11564 45444 11620 45726
rect 11228 44382 11230 44434
rect 11282 44382 11284 44434
rect 11228 44370 11284 44382
rect 11340 45388 11620 45444
rect 11676 45444 11732 45836
rect 11788 45668 11844 45678
rect 11788 45574 11844 45612
rect 11676 45388 11844 45444
rect 10556 43922 10612 43932
rect 10780 44044 11060 44100
rect 10668 43764 10724 43802
rect 10444 43652 10612 43708
rect 10668 43698 10724 43708
rect 9884 43598 9886 43650
rect 9938 43598 9940 43650
rect 9884 43586 9940 43598
rect 10444 43538 10500 43550
rect 10444 43486 10446 43538
rect 10498 43486 10500 43538
rect 9996 42868 10052 42878
rect 9996 42774 10052 42812
rect 9884 42756 9940 42766
rect 9884 42084 9940 42700
rect 10444 42532 10500 43486
rect 9884 41990 9940 42028
rect 9996 42308 10052 42318
rect 9996 42082 10052 42252
rect 10444 42196 10500 42476
rect 10556 42308 10612 43652
rect 10556 42242 10612 42252
rect 10668 43428 10724 43438
rect 10444 42130 10500 42140
rect 10668 42196 10724 43372
rect 10668 42130 10724 42140
rect 9996 42030 9998 42082
rect 10050 42030 10052 42082
rect 9996 42018 10052 42030
rect 10556 41972 10612 41982
rect 9772 41524 9828 41804
rect 10444 41970 10612 41972
rect 10444 41918 10558 41970
rect 10610 41918 10612 41970
rect 10444 41916 10612 41918
rect 9884 41748 9940 41758
rect 9884 41654 9940 41692
rect 9772 41468 10164 41524
rect 9996 41300 10052 41310
rect 9884 41298 10052 41300
rect 9884 41246 9998 41298
rect 10050 41246 10052 41298
rect 9884 41244 10052 41246
rect 9660 41188 9716 41198
rect 9884 41188 9940 41244
rect 9996 41234 10052 41244
rect 9660 40626 9716 41132
rect 9660 40574 9662 40626
rect 9714 40574 9716 40626
rect 9660 40404 9716 40574
rect 9660 40338 9716 40348
rect 9772 41132 9940 41188
rect 9772 39060 9828 41132
rect 9996 41076 10052 41086
rect 9884 40628 9940 40638
rect 9884 40514 9940 40572
rect 9884 40462 9886 40514
rect 9938 40462 9940 40514
rect 9996 40570 10052 41020
rect 9996 40518 9998 40570
rect 10050 40518 10052 40570
rect 9996 40506 10052 40518
rect 9884 40404 9940 40462
rect 10108 40404 10164 41468
rect 9884 40338 9940 40348
rect 9996 40348 10164 40404
rect 9996 40180 10052 40348
rect 9772 38994 9828 39004
rect 9884 40124 10052 40180
rect 9884 38162 9940 40124
rect 10108 39844 10164 39854
rect 10108 39618 10164 39788
rect 10108 39566 10110 39618
rect 10162 39566 10164 39618
rect 10108 39554 10164 39566
rect 10220 39396 10276 39406
rect 9884 38110 9886 38162
rect 9938 38110 9940 38162
rect 9884 38098 9940 38110
rect 9996 39172 10052 39182
rect 9996 38164 10052 39116
rect 10220 39058 10276 39340
rect 10220 39006 10222 39058
rect 10274 39006 10276 39058
rect 10220 38994 10276 39006
rect 10332 38948 10388 38958
rect 10220 38836 10276 38846
rect 10220 38742 10276 38780
rect 10332 38834 10388 38892
rect 10332 38782 10334 38834
rect 10386 38782 10388 38834
rect 10332 38724 10388 38782
rect 10332 38658 10388 38668
rect 9996 38098 10052 38108
rect 10332 37940 10388 37950
rect 10332 37846 10388 37884
rect 9996 37716 10052 37726
rect 10444 37716 10500 41916
rect 10556 41906 10612 41916
rect 10556 41300 10612 41310
rect 10556 40402 10612 41244
rect 10556 40350 10558 40402
rect 10610 40350 10612 40402
rect 10556 39844 10612 40350
rect 10780 40180 10836 44044
rect 11340 43988 11396 45388
rect 11452 45218 11508 45230
rect 11452 45166 11454 45218
rect 11506 45166 11508 45218
rect 11452 45108 11508 45166
rect 11452 45042 11508 45052
rect 11676 45108 11732 45118
rect 11452 44884 11508 44894
rect 11452 44546 11508 44828
rect 11452 44494 11454 44546
rect 11506 44494 11508 44546
rect 11452 44482 11508 44494
rect 10892 43932 11396 43988
rect 10892 43708 10948 43932
rect 11340 43764 11396 43774
rect 11564 43764 11620 43774
rect 10892 43652 11172 43708
rect 11340 43652 11508 43708
rect 10780 40124 11060 40180
rect 10556 39778 10612 39788
rect 10780 39508 10836 39518
rect 10780 39414 10836 39452
rect 10892 39396 10948 39406
rect 10556 39060 10612 39070
rect 10556 38834 10612 39004
rect 10556 38782 10558 38834
rect 10610 38782 10612 38834
rect 10556 38770 10612 38782
rect 10668 38164 10724 38174
rect 10668 38052 10724 38108
rect 9884 37492 9940 37502
rect 9548 35186 9604 35196
rect 9660 37044 9716 37054
rect 9436 34402 9492 34412
rect 9660 34356 9716 36988
rect 9884 37044 9940 37436
rect 9996 37490 10052 37660
rect 9996 37438 9998 37490
rect 10050 37438 10052 37490
rect 9996 37426 10052 37438
rect 10108 37660 10500 37716
rect 10556 38050 10724 38052
rect 10556 37998 10670 38050
rect 10722 37998 10724 38050
rect 10556 37996 10724 37998
rect 9884 36978 9940 36988
rect 10108 36820 10164 37660
rect 10108 36754 10164 36764
rect 10220 37492 10276 37502
rect 10220 36594 10276 37436
rect 10556 37380 10612 37996
rect 10668 37986 10724 37996
rect 10220 36542 10222 36594
rect 10274 36542 10276 36594
rect 10220 36530 10276 36542
rect 10332 37324 10612 37380
rect 9772 36372 9828 36382
rect 9772 36258 9828 36316
rect 9772 36206 9774 36258
rect 9826 36206 9828 36258
rect 9772 36148 9828 36206
rect 9772 36092 10052 36148
rect 9772 35812 9828 35822
rect 9772 35138 9828 35756
rect 9772 35086 9774 35138
rect 9826 35086 9828 35138
rect 9772 35026 9828 35086
rect 9772 34974 9774 35026
rect 9826 34974 9828 35026
rect 9772 34962 9828 34974
rect 9884 35586 9940 35598
rect 9884 35534 9886 35586
rect 9938 35534 9940 35586
rect 9884 34692 9940 35534
rect 9996 35588 10052 36092
rect 10220 35588 10276 35598
rect 9996 35532 10220 35588
rect 10220 35494 10276 35532
rect 10332 35308 10388 37324
rect 10444 37154 10500 37166
rect 10444 37102 10446 37154
rect 10498 37102 10500 37154
rect 10444 36036 10500 37102
rect 10556 37044 10612 37054
rect 10780 37044 10836 37054
rect 10556 36950 10612 36988
rect 10668 36988 10780 37044
rect 10668 36594 10724 36988
rect 10780 36978 10836 36988
rect 10668 36542 10670 36594
rect 10722 36542 10724 36594
rect 10668 36530 10724 36542
rect 10444 35970 10500 35980
rect 10780 35924 10836 35934
rect 10780 35830 10836 35868
rect 9884 34626 9940 34636
rect 10220 35252 10388 35308
rect 9772 34356 9828 34366
rect 9660 34354 9828 34356
rect 9660 34302 9774 34354
rect 9826 34302 9828 34354
rect 9660 34300 9828 34302
rect 9772 34290 9828 34300
rect 10220 34354 10276 35252
rect 10332 35140 10388 35150
rect 10332 35026 10388 35084
rect 10332 34974 10334 35026
rect 10386 34974 10388 35026
rect 10332 34962 10388 34974
rect 10220 34302 10222 34354
rect 10274 34302 10276 34354
rect 10220 34290 10276 34302
rect 10668 34692 10724 34702
rect 10556 34020 10612 34030
rect 10556 33926 10612 33964
rect 10668 30660 10724 34636
rect 10892 31780 10948 39340
rect 11004 38388 11060 40124
rect 11116 38500 11172 43652
rect 11452 43650 11508 43652
rect 11452 43598 11454 43650
rect 11506 43598 11508 43650
rect 11452 43586 11508 43598
rect 11228 43540 11284 43550
rect 11228 43446 11284 43484
rect 11452 42644 11508 42654
rect 11340 41858 11396 41870
rect 11340 41806 11342 41858
rect 11394 41806 11396 41858
rect 11340 41524 11396 41806
rect 11340 41458 11396 41468
rect 11340 40404 11396 40414
rect 11452 40404 11508 42588
rect 11340 40402 11508 40404
rect 11340 40350 11342 40402
rect 11394 40350 11508 40402
rect 11340 40348 11508 40350
rect 11340 40180 11396 40348
rect 11340 40114 11396 40124
rect 11116 38434 11172 38444
rect 11228 38722 11284 38734
rect 11452 38724 11508 38734
rect 11228 38670 11230 38722
rect 11282 38670 11284 38722
rect 11004 38322 11060 38332
rect 11228 38276 11284 38670
rect 11340 38722 11508 38724
rect 11340 38670 11454 38722
rect 11506 38670 11508 38722
rect 11340 38668 11508 38670
rect 11340 38388 11396 38668
rect 11452 38658 11508 38668
rect 11340 38322 11396 38332
rect 11452 38500 11508 38510
rect 11228 38164 11284 38220
rect 11452 38164 11508 38444
rect 11004 38108 11284 38164
rect 11340 38108 11508 38164
rect 11004 37268 11060 38108
rect 11116 37940 11172 37950
rect 11340 37940 11396 38108
rect 11564 38052 11620 43708
rect 11676 43762 11732 45052
rect 11788 44546 11844 45388
rect 11788 44494 11790 44546
rect 11842 44494 11844 44546
rect 11788 44482 11844 44494
rect 11676 43710 11678 43762
rect 11730 43710 11732 43762
rect 11676 43698 11732 43710
rect 11788 43988 11844 43998
rect 11788 43650 11844 43932
rect 11788 43598 11790 43650
rect 11842 43598 11844 43650
rect 11788 43586 11844 43598
rect 11676 43540 11732 43550
rect 11676 38668 11732 43484
rect 11788 40068 11844 40078
rect 11788 39058 11844 40012
rect 11788 39006 11790 39058
rect 11842 39006 11844 39058
rect 11788 38994 11844 39006
rect 11676 38612 11844 38668
rect 11172 37884 11284 37940
rect 11116 37874 11172 37884
rect 11228 37826 11284 37884
rect 11340 37874 11396 37884
rect 11452 37996 11620 38052
rect 11676 38500 11732 38510
rect 11228 37774 11230 37826
rect 11282 37774 11284 37826
rect 11228 37762 11284 37774
rect 11452 37490 11508 37996
rect 11452 37438 11454 37490
rect 11506 37438 11508 37490
rect 11452 37426 11508 37438
rect 11564 37826 11620 37838
rect 11564 37774 11566 37826
rect 11618 37774 11620 37826
rect 11004 36708 11060 37212
rect 11004 36642 11060 36652
rect 11116 37266 11172 37278
rect 11116 37214 11118 37266
rect 11170 37214 11172 37266
rect 11116 35700 11172 37214
rect 11228 36372 11284 36382
rect 11228 36278 11284 36316
rect 11004 34804 11060 34814
rect 11004 34468 11060 34748
rect 11004 34354 11060 34412
rect 11004 34302 11006 34354
rect 11058 34302 11060 34354
rect 11004 34290 11060 34302
rect 11004 33796 11060 33806
rect 11004 33458 11060 33740
rect 11116 33572 11172 35644
rect 11228 35588 11284 35598
rect 11228 35586 11396 35588
rect 11228 35534 11230 35586
rect 11282 35534 11396 35586
rect 11228 35532 11396 35534
rect 11228 35522 11284 35532
rect 11228 34916 11284 34926
rect 11228 34822 11284 34860
rect 11116 33506 11172 33516
rect 11004 33406 11006 33458
rect 11058 33406 11060 33458
rect 11004 33394 11060 33406
rect 10892 31714 10948 31724
rect 11340 31668 11396 35532
rect 11564 35140 11620 37774
rect 11676 36370 11732 38444
rect 11788 37044 11844 38612
rect 11788 36978 11844 36988
rect 11676 36318 11678 36370
rect 11730 36318 11732 36370
rect 11676 36260 11732 36318
rect 11676 36194 11732 36204
rect 11788 36148 11844 36158
rect 11676 35588 11732 35598
rect 11676 35494 11732 35532
rect 11564 35074 11620 35084
rect 11676 35138 11732 35150
rect 11676 35086 11678 35138
rect 11730 35086 11732 35138
rect 11564 34916 11620 34926
rect 11676 34916 11732 35086
rect 11564 34914 11732 34916
rect 11564 34862 11566 34914
rect 11618 34862 11732 34914
rect 11564 34860 11732 34862
rect 11564 34850 11620 34860
rect 11564 34580 11620 34590
rect 11564 34354 11620 34524
rect 11564 34302 11566 34354
rect 11618 34302 11620 34354
rect 11564 34290 11620 34302
rect 11340 31602 11396 31612
rect 11676 33460 11732 33470
rect 10668 30594 10724 30604
rect 9212 29698 9268 29708
rect 7756 24098 7812 24108
rect 7308 23202 7364 23212
rect 11676 21812 11732 33404
rect 11788 26908 11844 36092
rect 11900 32788 11956 45950
rect 12012 44882 12068 44894
rect 12012 44830 12014 44882
rect 12066 44830 12068 44882
rect 12012 43708 12068 44830
rect 12124 43988 12180 46956
rect 12236 46452 12292 49868
rect 21532 49924 21588 49934
rect 21532 49800 21588 49868
rect 32060 49924 32116 49934
rect 25788 49812 25844 49822
rect 26124 49812 26180 49822
rect 12768 49200 12880 49800
rect 14784 49200 14896 49800
rect 16128 49200 16240 49800
rect 17948 49588 18004 49598
rect 16828 49364 16884 49374
rect 12236 45330 12292 46396
rect 12348 47236 12404 47246
rect 12348 45668 12404 47180
rect 12684 46900 12740 46910
rect 12348 45602 12404 45612
rect 12460 45778 12516 45790
rect 12460 45726 12462 45778
rect 12514 45726 12516 45778
rect 12460 45444 12516 45726
rect 12460 45378 12516 45388
rect 12236 45278 12238 45330
rect 12290 45278 12292 45330
rect 12236 45266 12292 45278
rect 12348 44884 12404 44894
rect 12348 44790 12404 44828
rect 12124 43922 12180 43932
rect 12348 44660 12404 44670
rect 12348 44322 12404 44604
rect 12348 44270 12350 44322
rect 12402 44270 12404 44322
rect 12348 43764 12404 44270
rect 12572 44210 12628 44222
rect 12572 44158 12574 44210
rect 12626 44158 12628 44210
rect 12572 44100 12628 44158
rect 12572 44034 12628 44044
rect 12684 44098 12740 46844
rect 12796 46340 12852 49200
rect 15708 49140 15764 49150
rect 13804 49028 13860 49038
rect 13468 48020 13524 48030
rect 12796 46274 12852 46284
rect 13356 46452 13412 46462
rect 13356 46228 13412 46396
rect 13356 46162 13412 46172
rect 12796 45668 12852 45678
rect 12796 45666 13188 45668
rect 12796 45614 12798 45666
rect 12850 45614 13188 45666
rect 12796 45612 13188 45614
rect 12796 45602 12852 45612
rect 12908 44996 12964 45006
rect 12908 44902 12964 44940
rect 12908 44324 12964 44334
rect 12908 44230 12964 44268
rect 12684 44046 12686 44098
rect 12738 44046 12740 44098
rect 12684 44034 12740 44046
rect 12012 43652 12292 43708
rect 12348 43698 12404 43708
rect 13132 43708 13188 45612
rect 13244 45332 13300 45342
rect 13244 45106 13300 45276
rect 13244 45054 13246 45106
rect 13298 45054 13300 45106
rect 13244 45042 13300 45054
rect 13468 45218 13524 47964
rect 13580 45892 13636 45902
rect 13580 45798 13636 45836
rect 13468 45166 13470 45218
rect 13522 45166 13524 45218
rect 13468 44884 13524 45166
rect 13468 44818 13524 44828
rect 13692 44210 13748 44222
rect 13692 44158 13694 44210
rect 13746 44158 13748 44210
rect 13132 43652 13300 43708
rect 12012 42868 12068 42878
rect 12012 40852 12068 42812
rect 12236 42756 12292 43652
rect 13020 43540 13076 43550
rect 13020 43538 13188 43540
rect 13020 43486 13022 43538
rect 13074 43486 13188 43538
rect 13020 43484 13188 43486
rect 13020 43474 13076 43484
rect 12684 43426 12740 43438
rect 12684 43374 12686 43426
rect 12738 43374 12740 43426
rect 12684 43092 12740 43374
rect 12684 43026 12740 43036
rect 12236 42700 12628 42756
rect 12124 42644 12180 42654
rect 12124 42642 12404 42644
rect 12124 42590 12126 42642
rect 12178 42590 12404 42642
rect 12124 42588 12404 42590
rect 12124 42578 12180 42588
rect 12124 42196 12180 42206
rect 12124 41524 12180 42140
rect 12124 41076 12180 41468
rect 12124 41074 12292 41076
rect 12124 41022 12126 41074
rect 12178 41022 12292 41074
rect 12124 41020 12292 41022
rect 12124 41010 12180 41020
rect 12012 40796 12180 40852
rect 12124 38050 12180 40796
rect 12236 38500 12292 41020
rect 12236 38434 12292 38444
rect 12348 39844 12404 42588
rect 12348 38274 12404 39788
rect 12348 38222 12350 38274
rect 12402 38222 12404 38274
rect 12348 38210 12404 38222
rect 12460 39508 12516 39518
rect 12124 37998 12126 38050
rect 12178 37998 12180 38050
rect 12124 37986 12180 37998
rect 12460 38052 12516 39452
rect 12572 38500 12628 42700
rect 12908 42754 12964 42766
rect 12908 42702 12910 42754
rect 12962 42702 12964 42754
rect 12796 42308 12852 42318
rect 12572 38434 12628 38444
rect 12684 38724 12740 38734
rect 12684 38612 12740 38668
rect 12796 38668 12852 42252
rect 12908 41300 12964 42702
rect 13132 41748 13188 43484
rect 13132 41682 13188 41692
rect 12908 41186 12964 41244
rect 12908 41134 12910 41186
rect 12962 41134 12964 41186
rect 12908 41122 12964 41134
rect 12908 39844 12964 39854
rect 12908 39730 12964 39788
rect 12908 39678 12910 39730
rect 12962 39678 12964 39730
rect 12908 39666 12964 39678
rect 13244 39060 13300 43652
rect 13692 43652 13748 44158
rect 13804 44212 13860 48972
rect 14588 48804 14644 48814
rect 13916 47460 13972 47470
rect 13916 47366 13972 47404
rect 14140 47460 14196 47470
rect 14028 45108 14084 45118
rect 13804 44080 13860 44156
rect 13916 45052 14028 45108
rect 13916 43708 13972 45052
rect 14028 44976 14084 45052
rect 14028 44660 14084 44670
rect 14028 44322 14084 44604
rect 14028 44270 14030 44322
rect 14082 44270 14084 44322
rect 14028 44258 14084 44270
rect 13916 43652 14084 43708
rect 13692 43586 13748 43596
rect 13468 43540 13524 43550
rect 14028 43540 14084 43652
rect 13468 43538 13636 43540
rect 13468 43486 13470 43538
rect 13522 43486 13636 43538
rect 13468 43484 13636 43486
rect 13468 43474 13524 43484
rect 13468 41858 13524 41870
rect 13468 41806 13470 41858
rect 13522 41806 13524 41858
rect 13468 41748 13524 41806
rect 13468 40852 13524 41692
rect 13468 40786 13524 40796
rect 13468 40628 13524 40638
rect 13468 40290 13524 40572
rect 13580 40516 13636 43484
rect 14028 43446 14084 43484
rect 13692 43316 13748 43326
rect 13692 42754 13748 43260
rect 13692 42702 13694 42754
rect 13746 42702 13748 42754
rect 13692 42690 13748 42702
rect 14028 42756 14084 42766
rect 14140 42756 14196 47404
rect 14364 44772 14420 44782
rect 14364 43092 14420 44716
rect 14364 43026 14420 43036
rect 14476 44322 14532 44334
rect 14476 44270 14478 44322
rect 14530 44270 14532 44322
rect 14476 43540 14532 44270
rect 14028 42754 14196 42756
rect 14028 42702 14030 42754
rect 14082 42702 14196 42754
rect 14028 42700 14196 42702
rect 14476 42754 14532 43484
rect 14476 42702 14478 42754
rect 14530 42702 14532 42754
rect 14028 42690 14084 42700
rect 13804 42532 13860 42542
rect 13804 42530 13972 42532
rect 13804 42478 13806 42530
rect 13858 42478 13972 42530
rect 13804 42476 13972 42478
rect 13804 42466 13860 42476
rect 13916 42420 13972 42476
rect 13804 40964 13860 40974
rect 13580 40450 13636 40460
rect 13692 40908 13804 40964
rect 13468 40238 13470 40290
rect 13522 40238 13524 40290
rect 13468 40226 13524 40238
rect 13580 39508 13636 39518
rect 13580 39414 13636 39452
rect 13132 39004 13300 39060
rect 12908 38948 12964 38958
rect 12908 38834 12964 38892
rect 12908 38782 12910 38834
rect 12962 38782 12964 38834
rect 12908 38770 12964 38782
rect 13020 38836 13076 38846
rect 13020 38722 13076 38780
rect 13020 38670 13022 38722
rect 13074 38670 13076 38722
rect 12796 38612 12964 38668
rect 12572 38052 12628 38062
rect 12460 37996 12572 38052
rect 12572 37958 12628 37996
rect 12236 37828 12292 37838
rect 12124 37826 12292 37828
rect 12124 37774 12238 37826
rect 12290 37774 12292 37826
rect 12124 37772 12292 37774
rect 12124 37156 12180 37772
rect 12236 37762 12292 37772
rect 12236 37604 12292 37614
rect 12236 37490 12292 37548
rect 12236 37438 12238 37490
rect 12290 37438 12292 37490
rect 12236 37380 12292 37438
rect 12236 37314 12292 37324
rect 12348 37268 12404 37278
rect 12684 37268 12740 38556
rect 12124 37100 12292 37156
rect 12012 37042 12068 37054
rect 12012 36990 12014 37042
rect 12066 36990 12068 37042
rect 12012 36932 12068 36990
rect 12012 36866 12068 36876
rect 12012 36260 12068 36270
rect 12012 36166 12068 36204
rect 12012 35586 12068 35598
rect 12012 35534 12014 35586
rect 12066 35534 12068 35586
rect 12012 35476 12068 35534
rect 12012 35138 12068 35420
rect 12012 35086 12014 35138
rect 12066 35086 12068 35138
rect 12012 35026 12068 35086
rect 12012 34974 12014 35026
rect 12066 34974 12068 35026
rect 12012 34962 12068 34974
rect 12124 34580 12180 34590
rect 12012 34356 12068 34366
rect 12124 34356 12180 34524
rect 12012 34354 12180 34356
rect 12012 34302 12014 34354
rect 12066 34302 12180 34354
rect 12012 34300 12180 34302
rect 12012 34290 12068 34300
rect 12124 33460 12180 33470
rect 12124 33366 12180 33404
rect 11900 32722 11956 32732
rect 12236 32676 12292 37100
rect 12348 37154 12404 37212
rect 12348 37102 12350 37154
rect 12402 37102 12404 37154
rect 12348 37090 12404 37102
rect 12460 37212 12740 37268
rect 12796 38050 12852 38062
rect 12796 37998 12798 38050
rect 12850 37998 12852 38050
rect 12348 36260 12404 36270
rect 12348 33348 12404 36204
rect 12460 35812 12516 37212
rect 12796 37156 12852 37998
rect 12572 37100 12852 37156
rect 12572 36820 12628 37100
rect 12908 37044 12964 38612
rect 12572 36484 12628 36764
rect 12572 36418 12628 36428
rect 12796 37042 12964 37044
rect 12796 36990 12910 37042
rect 12962 36990 12964 37042
rect 12796 36988 12964 36990
rect 12572 36258 12628 36270
rect 12572 36206 12574 36258
rect 12626 36206 12628 36258
rect 12572 36148 12628 36206
rect 12572 36082 12628 36092
rect 12572 35812 12628 35822
rect 12516 35810 12628 35812
rect 12516 35758 12574 35810
rect 12626 35758 12628 35810
rect 12516 35756 12628 35758
rect 12460 35680 12516 35756
rect 12572 35746 12628 35756
rect 12684 35474 12740 35486
rect 12684 35422 12686 35474
rect 12738 35422 12740 35474
rect 12684 34916 12740 35422
rect 12684 34850 12740 34860
rect 12572 34692 12628 34702
rect 12628 34636 12740 34692
rect 12572 34560 12628 34636
rect 12460 34356 12516 34366
rect 12460 33908 12516 34300
rect 12460 33842 12516 33852
rect 12572 33684 12628 33694
rect 12572 33458 12628 33628
rect 12572 33406 12574 33458
rect 12626 33406 12628 33458
rect 12572 33394 12628 33406
rect 12348 33282 12404 33292
rect 12236 32610 12292 32620
rect 12572 33236 12628 33246
rect 12572 32786 12628 33180
rect 12572 32734 12574 32786
rect 12626 32734 12628 32786
rect 12236 32452 12292 32462
rect 12236 32358 12292 32396
rect 12572 32004 12628 32734
rect 12572 31938 12628 31948
rect 12684 26908 12740 34636
rect 12796 33796 12852 36988
rect 12908 36978 12964 36988
rect 12908 36370 12964 36382
rect 12908 36318 12910 36370
rect 12962 36318 12964 36370
rect 12908 36260 12964 36318
rect 12908 36194 12964 36204
rect 13020 36148 13076 38670
rect 13020 36082 13076 36092
rect 12908 36036 12964 36046
rect 12908 34354 12964 35980
rect 13132 36036 13188 39004
rect 13356 38724 13412 38734
rect 13356 38630 13412 38668
rect 13692 38276 13748 40908
rect 13804 40870 13860 40908
rect 13916 40292 13972 42364
rect 14140 41972 14196 41982
rect 14476 41972 14532 42702
rect 14588 43652 14644 48748
rect 14812 48804 14868 48814
rect 14812 48468 14868 48748
rect 14812 48402 14868 48412
rect 14700 47684 14756 47694
rect 14700 47234 14756 47628
rect 14700 47182 14702 47234
rect 14754 47182 14756 47234
rect 14700 47170 14756 47182
rect 15484 47458 15540 47470
rect 15484 47406 15486 47458
rect 15538 47406 15540 47458
rect 15260 46676 15316 46686
rect 15260 45444 15316 46620
rect 15148 45332 15204 45342
rect 14588 42084 14644 43596
rect 14588 42018 14644 42028
rect 14700 45220 14756 45230
rect 14140 41970 14532 41972
rect 14140 41918 14142 41970
rect 14194 41918 14532 41970
rect 14140 41916 14532 41918
rect 14140 41300 14196 41916
rect 14028 41076 14084 41086
rect 14028 40982 14084 41020
rect 13916 40226 13972 40236
rect 14140 40402 14196 41244
rect 14476 41300 14532 41310
rect 14476 41206 14532 41244
rect 14588 41188 14644 41198
rect 14588 41094 14644 41132
rect 14140 40350 14142 40402
rect 14194 40350 14196 40402
rect 13916 39620 13972 39630
rect 13916 39506 13972 39564
rect 13916 39454 13918 39506
rect 13970 39454 13972 39506
rect 13804 39394 13860 39406
rect 13804 39342 13806 39394
rect 13858 39342 13860 39394
rect 13804 39284 13860 39342
rect 13804 39218 13860 39228
rect 13916 38836 13972 39454
rect 13916 38770 13972 38780
rect 14028 39060 14084 39070
rect 14028 38668 14084 39004
rect 13692 38210 13748 38220
rect 13916 38612 14084 38668
rect 14140 38834 14196 40350
rect 14476 39730 14532 39742
rect 14476 39678 14478 39730
rect 14530 39678 14532 39730
rect 14476 39620 14532 39678
rect 14476 39554 14532 39564
rect 14700 38948 14756 45164
rect 14812 44996 14868 45006
rect 14812 44994 15092 44996
rect 14812 44942 14814 44994
rect 14866 44942 15092 44994
rect 14812 44940 15092 44942
rect 14812 44930 14868 44940
rect 14812 43652 14868 43662
rect 14812 43558 14868 43596
rect 15036 42868 15092 44940
rect 15036 42802 15092 42812
rect 15148 43764 15204 45276
rect 15260 44434 15316 45388
rect 15260 44382 15262 44434
rect 15314 44382 15316 44434
rect 15260 44370 15316 44382
rect 15372 45778 15428 45790
rect 15372 45726 15374 45778
rect 15426 45726 15428 45778
rect 15372 45108 15428 45726
rect 15372 44324 15428 45052
rect 15372 44258 15428 44268
rect 15484 43708 15540 47406
rect 14812 42420 14868 42430
rect 14812 41970 14868 42364
rect 14812 41918 14814 41970
rect 14866 41918 14868 41970
rect 14812 41906 14868 41918
rect 15148 41300 15204 43708
rect 15260 43652 15540 43708
rect 15708 43988 15764 49084
rect 16828 49028 16884 49308
rect 16828 48962 16884 48972
rect 16492 48692 16548 48702
rect 15260 42866 15316 43652
rect 15260 42814 15262 42866
rect 15314 42814 15316 42866
rect 15260 42802 15316 42814
rect 15596 42084 15652 42094
rect 15148 41234 15204 41244
rect 15260 41412 15316 41422
rect 15260 41186 15316 41356
rect 15260 41134 15262 41186
rect 15314 41134 15316 41186
rect 15260 41122 15316 41134
rect 15596 41186 15652 42028
rect 15596 41134 15598 41186
rect 15650 41134 15652 41186
rect 14812 40404 14868 40414
rect 15596 40404 15652 41134
rect 14812 40310 14868 40348
rect 15036 40348 15652 40404
rect 14812 38948 14868 38958
rect 14700 38946 14868 38948
rect 14700 38894 14814 38946
rect 14866 38894 14868 38946
rect 14700 38892 14868 38894
rect 14812 38882 14868 38892
rect 14140 38782 14142 38834
rect 14194 38782 14196 38834
rect 14140 38668 14196 38782
rect 15036 38724 15092 40348
rect 15708 39620 15764 43932
rect 15820 47908 15876 47918
rect 15820 47236 15876 47852
rect 15820 43708 15876 47180
rect 16044 47236 16100 47246
rect 16044 47142 16100 47180
rect 16044 44212 16100 44222
rect 15820 43652 15988 43708
rect 14700 38668 15092 38724
rect 15484 39564 15764 39620
rect 15820 41412 15876 41422
rect 14140 38612 14644 38668
rect 13692 37940 13748 37950
rect 13692 37846 13748 37884
rect 13804 37826 13860 37838
rect 13804 37774 13806 37826
rect 13858 37774 13860 37826
rect 13804 37604 13860 37774
rect 13804 37538 13860 37548
rect 13468 37266 13524 37278
rect 13468 37214 13470 37266
rect 13522 37214 13524 37266
rect 13468 37156 13524 37214
rect 13916 37156 13972 38612
rect 14364 38500 14420 38510
rect 14028 38164 14084 38174
rect 14028 38050 14084 38108
rect 14028 37998 14030 38050
rect 14082 37998 14084 38050
rect 14028 37986 14084 37998
rect 14140 37940 14196 37950
rect 13468 37090 13524 37100
rect 13804 37100 13972 37156
rect 14028 37380 14084 37390
rect 14028 37154 14084 37324
rect 14028 37102 14030 37154
rect 14082 37102 14084 37154
rect 13244 37042 13300 37054
rect 13804 37044 13860 37100
rect 13244 36990 13246 37042
rect 13298 36990 13300 37042
rect 13244 36260 13300 36990
rect 13580 36988 13860 37044
rect 13244 36194 13300 36204
rect 13356 36820 13412 36830
rect 13132 35970 13188 35980
rect 13244 35700 13300 35710
rect 13132 35698 13300 35700
rect 13132 35646 13246 35698
rect 13298 35646 13300 35698
rect 13132 35644 13300 35646
rect 12908 34302 12910 34354
rect 12962 34302 12964 34354
rect 12908 34290 12964 34302
rect 13020 34690 13076 34702
rect 13020 34638 13022 34690
rect 13074 34638 13076 34690
rect 12796 33730 12852 33740
rect 13020 33348 13076 34638
rect 13020 33282 13076 33292
rect 13020 33122 13076 33134
rect 13020 33070 13022 33122
rect 13074 33070 13076 33122
rect 13020 33012 13076 33070
rect 13020 32946 13076 32956
rect 13132 32450 13188 35644
rect 13244 35634 13300 35644
rect 13244 34132 13300 34142
rect 13244 34038 13300 34076
rect 13356 33348 13412 36764
rect 13580 35922 13636 36988
rect 14028 36708 14084 37102
rect 13916 36652 14084 36708
rect 13804 36596 13860 36606
rect 13692 36370 13748 36382
rect 13692 36318 13694 36370
rect 13746 36318 13748 36370
rect 13692 36148 13748 36318
rect 13804 36370 13860 36540
rect 13804 36318 13806 36370
rect 13858 36318 13860 36370
rect 13804 36260 13860 36318
rect 13804 36194 13860 36204
rect 13692 36082 13748 36092
rect 13580 35870 13582 35922
rect 13634 35870 13636 35922
rect 13580 35858 13636 35870
rect 13468 35700 13524 35710
rect 13468 34468 13524 35644
rect 13916 35588 13972 36652
rect 14028 36484 14084 36494
rect 14028 36390 14084 36428
rect 14140 35812 14196 37884
rect 13468 34402 13524 34412
rect 13580 35532 13972 35588
rect 14028 35810 14196 35812
rect 14028 35758 14142 35810
rect 14194 35758 14196 35810
rect 14028 35756 14196 35758
rect 13580 33460 13636 35532
rect 13804 35252 13860 35262
rect 13804 35140 13860 35196
rect 13804 35084 13972 35140
rect 13804 34804 13860 34814
rect 13692 34468 13748 34478
rect 13692 34354 13748 34412
rect 13692 34302 13694 34354
rect 13746 34302 13748 34354
rect 13692 34290 13748 34302
rect 13580 33394 13636 33404
rect 13692 33570 13748 33582
rect 13692 33518 13694 33570
rect 13746 33518 13748 33570
rect 13356 33282 13412 33292
rect 13580 33122 13636 33134
rect 13580 33070 13582 33122
rect 13634 33070 13636 33122
rect 13580 32900 13636 33070
rect 13580 32834 13636 32844
rect 13580 32676 13636 32686
rect 13692 32676 13748 33518
rect 13580 32674 13748 32676
rect 13580 32622 13582 32674
rect 13634 32622 13748 32674
rect 13580 32620 13748 32622
rect 13580 32610 13636 32620
rect 13132 32398 13134 32450
rect 13186 32398 13188 32450
rect 11788 26852 12404 26908
rect 12684 26852 12964 26908
rect 12348 26292 12404 26852
rect 12348 26226 12404 26236
rect 12908 23716 12964 26852
rect 13132 24948 13188 32398
rect 13804 31444 13860 34748
rect 13804 31378 13860 31388
rect 13916 29876 13972 35084
rect 14028 32900 14084 35756
rect 14140 35746 14196 35756
rect 14252 36932 14308 36942
rect 14140 34804 14196 34814
rect 14252 34804 14308 36876
rect 14364 35924 14420 38444
rect 14588 38050 14644 38612
rect 14588 37998 14590 38050
rect 14642 37998 14644 38050
rect 14588 36596 14644 37998
rect 14588 36482 14644 36540
rect 14588 36430 14590 36482
rect 14642 36430 14644 36482
rect 14476 35924 14532 35934
rect 14364 35868 14476 35924
rect 14476 35792 14532 35868
rect 14588 35700 14644 36430
rect 14140 34802 14308 34804
rect 14140 34750 14142 34802
rect 14194 34750 14308 34802
rect 14140 34748 14308 34750
rect 14364 35644 14644 35700
rect 14364 35476 14420 35644
rect 14140 34738 14196 34748
rect 14364 34580 14420 35420
rect 14700 34804 14756 38668
rect 15260 37940 15316 37950
rect 15148 37938 15316 37940
rect 15148 37886 15262 37938
rect 15314 37886 15316 37938
rect 15148 37884 15316 37886
rect 14700 34710 14756 34748
rect 14812 37604 14868 37614
rect 14140 34524 14420 34580
rect 14140 34018 14196 34524
rect 14140 33966 14142 34018
rect 14194 33966 14196 34018
rect 14140 33458 14196 33966
rect 14140 33406 14142 33458
rect 14194 33406 14196 33458
rect 14140 33394 14196 33406
rect 14252 34356 14308 34366
rect 14028 32844 14196 32900
rect 14028 32452 14084 32462
rect 14028 32358 14084 32396
rect 14140 31220 14196 32844
rect 14252 31890 14308 34300
rect 14700 34130 14756 34142
rect 14700 34078 14702 34130
rect 14754 34078 14756 34130
rect 14700 33684 14756 34078
rect 14812 34020 14868 37548
rect 15036 36148 15092 36158
rect 15036 35700 15092 36092
rect 15036 35606 15092 35644
rect 14924 35252 14980 35262
rect 14924 35026 14980 35196
rect 14924 34974 14926 35026
rect 14978 34974 14980 35026
rect 14924 34962 14980 34974
rect 14924 34690 14980 34702
rect 14924 34638 14926 34690
rect 14978 34638 14980 34690
rect 14924 34356 14980 34638
rect 14924 34290 14980 34300
rect 15036 34356 15092 34366
rect 15148 34356 15204 37884
rect 15260 37874 15316 37884
rect 15260 37268 15316 37278
rect 15260 36594 15316 37212
rect 15260 36542 15262 36594
rect 15314 36542 15316 36594
rect 15260 36530 15316 36542
rect 15372 36708 15428 36718
rect 15372 35698 15428 36652
rect 15484 35922 15540 39564
rect 15484 35870 15486 35922
rect 15538 35870 15540 35922
rect 15484 35858 15540 35870
rect 15708 35924 15764 35934
rect 15820 35924 15876 41356
rect 15932 38668 15988 43652
rect 16044 41076 16100 44156
rect 16492 41188 16548 48636
rect 16940 48468 16996 48478
rect 16940 47796 16996 48412
rect 16940 47730 16996 47740
rect 17836 47796 17892 47806
rect 16940 47572 16996 47582
rect 16716 47516 16940 47572
rect 16716 47458 16772 47516
rect 16940 47506 16996 47516
rect 16716 47406 16718 47458
rect 16770 47406 16772 47458
rect 16716 47394 16772 47406
rect 17388 46004 17444 46014
rect 16492 41122 16548 41132
rect 16604 45892 16660 45902
rect 16604 45444 16660 45836
rect 16044 41074 16436 41076
rect 16044 41022 16046 41074
rect 16098 41022 16436 41074
rect 16044 41020 16436 41022
rect 16044 41010 16100 41020
rect 15932 38612 16212 38668
rect 16156 38276 16212 38612
rect 16156 37378 16212 38220
rect 16156 37326 16158 37378
rect 16210 37326 16212 37378
rect 16156 37314 16212 37326
rect 15820 35868 16212 35924
rect 15372 35646 15374 35698
rect 15426 35646 15428 35698
rect 15372 35634 15428 35646
rect 15596 35700 15652 35710
rect 15596 35606 15652 35644
rect 15596 35364 15652 35374
rect 15708 35364 15764 35868
rect 15652 35308 15764 35364
rect 16044 35700 16100 35710
rect 15596 34804 15652 35308
rect 15820 35140 15876 35150
rect 15036 34354 15204 34356
rect 15036 34302 15038 34354
rect 15090 34302 15204 34354
rect 15036 34300 15204 34302
rect 15372 34802 15652 34804
rect 15372 34750 15598 34802
rect 15650 34750 15652 34802
rect 15372 34748 15652 34750
rect 15036 34290 15092 34300
rect 15372 34132 15428 34748
rect 15596 34738 15652 34748
rect 15708 35026 15764 35038
rect 15708 34974 15710 35026
rect 15762 34974 15764 35026
rect 15036 34076 15428 34132
rect 15596 34130 15652 34142
rect 15596 34078 15598 34130
rect 15650 34078 15652 34130
rect 14924 34020 14980 34030
rect 14812 33964 14924 34020
rect 14700 33618 14756 33628
rect 14588 33236 14644 33246
rect 14588 33142 14644 33180
rect 14924 33124 14980 33964
rect 15036 33570 15092 34076
rect 15596 34020 15652 34078
rect 15036 33518 15038 33570
rect 15090 33518 15092 33570
rect 15036 33506 15092 33518
rect 15148 33964 15652 34020
rect 15036 33348 15092 33358
rect 15036 33254 15092 33292
rect 14924 33068 15092 33124
rect 14924 32788 14980 32798
rect 14924 32694 14980 32732
rect 14476 32450 14532 32462
rect 14476 32398 14478 32450
rect 14530 32398 14532 32450
rect 14476 32340 14532 32398
rect 14476 32274 14532 32284
rect 14252 31838 14254 31890
rect 14306 31838 14308 31890
rect 14252 31826 14308 31838
rect 14700 31556 14756 31566
rect 14700 31462 14756 31500
rect 14140 31154 14196 31164
rect 14812 31220 14868 31230
rect 14812 30772 14868 31164
rect 15036 31220 15092 33068
rect 15036 31154 15092 31164
rect 15148 31554 15204 33964
rect 15708 33908 15764 34974
rect 15820 34914 15876 35084
rect 15820 34862 15822 34914
rect 15874 34862 15876 34914
rect 15820 34850 15876 34862
rect 16044 34802 16100 35644
rect 16044 34750 16046 34802
rect 16098 34750 16100 34802
rect 15932 34692 15988 34702
rect 15484 33852 15764 33908
rect 15820 34580 15876 34590
rect 15484 33684 15540 33852
rect 15820 33796 15876 34524
rect 15932 34354 15988 34636
rect 15932 34302 15934 34354
rect 15986 34302 15988 34354
rect 15932 34244 15988 34302
rect 15932 34178 15988 34188
rect 15372 33628 15540 33684
rect 15596 33740 15876 33796
rect 15372 32788 15428 33628
rect 15484 33460 15540 33470
rect 15484 33366 15540 33404
rect 15596 33236 15652 33740
rect 15148 31502 15150 31554
rect 15202 31502 15204 31554
rect 14812 30706 14868 30716
rect 15148 29988 15204 31502
rect 15148 29922 15204 29932
rect 15260 32732 15428 32788
rect 15484 33180 15652 33236
rect 15820 33572 15876 33582
rect 15820 33458 15876 33516
rect 15820 33406 15822 33458
rect 15874 33406 15876 33458
rect 15260 30100 15316 32732
rect 15372 32564 15428 32574
rect 15372 32470 15428 32508
rect 13916 29810 13972 29820
rect 15260 28644 15316 30044
rect 13132 24882 13188 24892
rect 15036 28588 15316 28644
rect 12908 23650 12964 23660
rect 11676 21746 11732 21756
rect 15036 16436 15092 28588
rect 15484 27524 15540 33180
rect 15820 33124 15876 33406
rect 15820 33058 15876 33068
rect 15596 32676 15652 32686
rect 16044 32676 16100 34750
rect 16156 35698 16212 35868
rect 16380 35700 16436 41020
rect 16492 39844 16548 39854
rect 16492 39508 16548 39788
rect 16604 39732 16660 45388
rect 16716 45666 16772 45678
rect 16716 45614 16718 45666
rect 16770 45614 16772 45666
rect 16716 45108 16772 45614
rect 17388 45108 17444 45948
rect 17724 46004 17780 46014
rect 17724 45910 17780 45948
rect 17724 45108 17780 45118
rect 17388 45052 17556 45108
rect 16716 41860 16772 45052
rect 16940 44996 16996 45006
rect 16940 44994 17108 44996
rect 16940 44942 16942 44994
rect 16994 44942 17108 44994
rect 16940 44940 17108 44942
rect 16940 44930 16996 44940
rect 17052 43540 17108 44940
rect 16940 43426 16996 43438
rect 16940 43374 16942 43426
rect 16994 43374 16996 43426
rect 16940 43316 16996 43374
rect 16940 43250 16996 43260
rect 17052 42644 17108 43484
rect 17388 44434 17444 44446
rect 17388 44382 17390 44434
rect 17442 44382 17444 44434
rect 17052 42578 17108 42588
rect 17276 43428 17332 43438
rect 16716 41794 16772 41804
rect 16940 42084 16996 42094
rect 16940 41858 16996 42028
rect 16940 41806 16942 41858
rect 16994 41806 16996 41858
rect 16940 41794 16996 41806
rect 17052 41524 17108 41534
rect 17052 41186 17108 41468
rect 17052 41134 17054 41186
rect 17106 41134 17108 41186
rect 17052 41122 17108 41134
rect 16716 41074 16772 41086
rect 16716 41022 16718 41074
rect 16770 41022 16772 41074
rect 16716 40852 16772 41022
rect 17276 41076 17332 43372
rect 17388 43204 17444 44382
rect 17388 43138 17444 43148
rect 17388 42868 17444 42878
rect 17388 42774 17444 42812
rect 17500 42308 17556 45052
rect 17724 45014 17780 45052
rect 17836 44884 17892 47740
rect 17612 44828 17892 44884
rect 17612 43428 17668 44828
rect 17948 44772 18004 49532
rect 18144 49200 18256 49800
rect 20160 49200 20272 49800
rect 21504 49200 21616 49800
rect 23212 49364 23268 49374
rect 17836 44716 18004 44772
rect 18060 49140 18116 49150
rect 17612 43362 17668 43372
rect 17724 44324 17780 44334
rect 17724 42756 17780 44268
rect 17836 43652 17892 44716
rect 17948 44324 18004 44334
rect 17948 44230 18004 44268
rect 17836 43586 17892 43596
rect 17948 43650 18004 43662
rect 17948 43598 17950 43650
rect 18002 43598 18004 43650
rect 17948 43428 18004 43598
rect 17948 43362 18004 43372
rect 17948 42756 18004 42766
rect 17724 42754 18004 42756
rect 17724 42702 17950 42754
rect 18002 42702 18004 42754
rect 17724 42700 18004 42702
rect 17948 42690 18004 42700
rect 17500 42252 18004 42308
rect 17836 42084 17892 42094
rect 17836 41970 17892 42028
rect 17836 41918 17838 41970
rect 17890 41918 17892 41970
rect 17836 41906 17892 41918
rect 17948 41746 18004 42252
rect 18060 42196 18116 49084
rect 18172 45780 18228 49200
rect 18172 45714 18228 45724
rect 18284 49028 18340 49038
rect 18284 43708 18340 48972
rect 18956 48692 19012 48702
rect 18060 42130 18116 42140
rect 18172 43652 18340 43708
rect 18508 47348 18564 47358
rect 18396 43652 18452 43662
rect 18172 41972 18228 43652
rect 18172 41906 18228 41916
rect 18284 42194 18340 42206
rect 18284 42142 18286 42194
rect 18338 42142 18340 42194
rect 18172 41748 18228 41758
rect 17948 41694 17950 41746
rect 18002 41694 18004 41746
rect 17276 41010 17332 41020
rect 17388 41300 17444 41310
rect 16716 40786 16772 40796
rect 16940 40292 16996 40302
rect 16940 40290 17108 40292
rect 16940 40238 16942 40290
rect 16994 40238 17108 40290
rect 16940 40236 17108 40238
rect 16940 40226 16996 40236
rect 16604 39676 16772 39732
rect 16604 39508 16660 39518
rect 16492 39506 16660 39508
rect 16492 39454 16606 39506
rect 16658 39454 16660 39506
rect 16492 39452 16660 39454
rect 16156 35646 16158 35698
rect 16210 35646 16212 35698
rect 16156 34580 16212 35646
rect 16268 35698 16436 35700
rect 16268 35646 16382 35698
rect 16434 35646 16436 35698
rect 16268 35644 16436 35646
rect 16268 34804 16324 35644
rect 16380 35634 16436 35644
rect 16492 38164 16548 38174
rect 16492 35476 16548 38108
rect 16604 37044 16660 39452
rect 16604 36978 16660 36988
rect 16604 35924 16660 35934
rect 16604 35830 16660 35868
rect 16268 34738 16324 34748
rect 16380 35420 16548 35476
rect 16604 35476 16660 35486
rect 16156 34514 16212 34524
rect 16380 34580 16436 35420
rect 16604 35382 16660 35420
rect 16492 35140 16548 35150
rect 16492 35046 16548 35084
rect 16380 34514 16436 34524
rect 16716 34468 16772 39676
rect 16940 38722 16996 38734
rect 16940 38670 16942 38722
rect 16994 38670 16996 38722
rect 16828 37266 16884 37278
rect 16828 37214 16830 37266
rect 16882 37214 16884 37266
rect 16828 36596 16884 37214
rect 16828 36530 16884 36540
rect 16940 35924 16996 38670
rect 17052 38388 17108 40236
rect 17052 38322 17108 38332
rect 17276 39618 17332 39630
rect 17276 39566 17278 39618
rect 17330 39566 17332 39618
rect 17276 37940 17332 39566
rect 17388 38164 17444 41244
rect 17500 41188 17556 41198
rect 17500 41094 17556 41132
rect 17836 40964 17892 40974
rect 17724 40962 17892 40964
rect 17724 40910 17838 40962
rect 17890 40910 17892 40962
rect 17724 40908 17892 40910
rect 17612 40740 17668 40750
rect 17612 40402 17668 40684
rect 17612 40350 17614 40402
rect 17666 40350 17668 40402
rect 17612 40338 17668 40350
rect 17388 38070 17444 38108
rect 17612 38722 17668 38734
rect 17612 38670 17614 38722
rect 17666 38670 17668 38722
rect 17612 38610 17668 38670
rect 17612 38558 17614 38610
rect 17666 38558 17668 38610
rect 17612 37940 17668 38558
rect 17276 37884 17668 37940
rect 17276 36596 17332 37884
rect 17276 36530 17332 36540
rect 17388 36820 17444 36830
rect 17612 36820 17668 36830
rect 17388 36594 17444 36764
rect 17388 36542 17390 36594
rect 17442 36542 17444 36594
rect 16940 35868 17332 35924
rect 16940 35700 16996 35710
rect 16940 35606 16996 35644
rect 16716 34402 16772 34412
rect 16940 34914 16996 34926
rect 16940 34862 16942 34914
rect 16994 34862 16996 34914
rect 16492 34244 16548 34254
rect 16380 34242 16548 34244
rect 16380 34190 16494 34242
rect 16546 34190 16548 34242
rect 16380 34188 16548 34190
rect 16380 33572 16436 34188
rect 16492 34178 16548 34188
rect 16716 34132 16772 34142
rect 16716 34038 16772 34076
rect 16604 34020 16660 34030
rect 16604 33926 16660 33964
rect 16380 33516 16548 33572
rect 16268 33124 16324 33134
rect 15596 31890 15652 32620
rect 15820 32620 16100 32676
rect 16156 33012 16212 33022
rect 16156 32786 16212 32956
rect 16156 32734 16158 32786
rect 16210 32734 16212 32786
rect 15708 32450 15764 32462
rect 15708 32398 15710 32450
rect 15762 32398 15764 32450
rect 15708 32116 15764 32398
rect 15708 32050 15764 32060
rect 15596 31838 15598 31890
rect 15650 31838 15652 31890
rect 15596 31826 15652 31838
rect 15596 30996 15652 31006
rect 15596 30902 15652 30940
rect 15820 30660 15876 32620
rect 16156 32228 16212 32734
rect 16044 31668 16100 31678
rect 16044 31574 16100 31612
rect 16156 31108 16212 32172
rect 15820 30594 15876 30604
rect 16044 31052 16212 31108
rect 16268 32004 16324 33068
rect 16380 33122 16436 33134
rect 16380 33070 16382 33122
rect 16434 33070 16436 33122
rect 16380 33012 16436 33070
rect 16380 32946 16436 32956
rect 16044 30212 16100 31052
rect 16156 30882 16212 30894
rect 16156 30830 16158 30882
rect 16210 30830 16212 30882
rect 16156 30770 16212 30830
rect 16156 30718 16158 30770
rect 16210 30718 16212 30770
rect 16156 30706 16212 30718
rect 16044 30146 16100 30156
rect 16156 30212 16212 30222
rect 16268 30212 16324 31948
rect 16380 31780 16436 31790
rect 16380 31332 16436 31724
rect 16380 31266 16436 31276
rect 16492 30770 16548 33516
rect 16716 33122 16772 33134
rect 16716 33070 16718 33122
rect 16770 33070 16772 33122
rect 16716 33012 16772 33070
rect 16716 32946 16772 32956
rect 16828 32788 16884 32798
rect 16828 32694 16884 32732
rect 16716 32676 16772 32686
rect 16716 32582 16772 32620
rect 16828 32340 16884 32350
rect 16940 32340 16996 34862
rect 17164 34914 17220 34926
rect 17164 34862 17166 34914
rect 17218 34862 17220 34914
rect 17052 34130 17108 34142
rect 17052 34078 17054 34130
rect 17106 34078 17108 34130
rect 17052 33796 17108 34078
rect 17052 33730 17108 33740
rect 17052 33348 17108 33358
rect 17052 32786 17108 33292
rect 17052 32734 17054 32786
rect 17106 32734 17108 32786
rect 17052 32722 17108 32734
rect 16884 32284 16996 32340
rect 17052 32340 17108 32350
rect 16716 31892 16772 31902
rect 16604 31220 16660 31230
rect 16716 31220 16772 31836
rect 16604 31218 16772 31220
rect 16604 31166 16606 31218
rect 16658 31166 16772 31218
rect 16604 31164 16772 31166
rect 16604 31154 16660 31164
rect 16492 30718 16494 30770
rect 16546 30718 16548 30770
rect 16492 30706 16548 30718
rect 16716 30770 16772 30782
rect 16716 30718 16718 30770
rect 16770 30718 16772 30770
rect 16156 30210 16324 30212
rect 16156 30158 16158 30210
rect 16210 30158 16324 30210
rect 16156 30156 16324 30158
rect 16604 30660 16660 30670
rect 15484 27458 15540 27468
rect 16156 16772 16212 30156
rect 16604 29316 16660 30604
rect 16604 29250 16660 29260
rect 16716 26404 16772 30718
rect 16828 30660 16884 32284
rect 16940 31554 16996 31566
rect 16940 31502 16942 31554
rect 16994 31502 16996 31554
rect 16940 31444 16996 31502
rect 16940 31220 16996 31388
rect 16940 31154 16996 31164
rect 17052 31218 17108 32284
rect 17052 31166 17054 31218
rect 17106 31166 17108 31218
rect 17052 31154 17108 31166
rect 16828 30594 16884 30604
rect 17164 30996 17220 34862
rect 17276 33572 17332 35868
rect 17388 35252 17444 36542
rect 17388 35186 17444 35196
rect 17500 36764 17612 36820
rect 17500 35476 17556 36764
rect 17612 36754 17668 36764
rect 17724 36260 17780 40908
rect 17836 40898 17892 40908
rect 17948 40740 18004 41694
rect 17836 40684 18004 40740
rect 18060 41746 18228 41748
rect 18060 41694 18174 41746
rect 18226 41694 18228 41746
rect 18060 41692 18228 41694
rect 17836 39620 17892 40684
rect 18060 40628 18116 41692
rect 18172 41682 18228 41692
rect 17948 40572 18116 40628
rect 18172 41076 18228 41086
rect 18172 40626 18228 41020
rect 18172 40574 18174 40626
rect 18226 40574 18228 40626
rect 17948 39844 18004 40572
rect 18172 40562 18228 40574
rect 18284 40628 18340 42142
rect 18396 42196 18452 43596
rect 18508 43540 18564 47292
rect 18732 47124 18788 47134
rect 18620 45220 18676 45230
rect 18620 45126 18676 45164
rect 18732 44434 18788 47068
rect 18732 44382 18734 44434
rect 18786 44382 18788 44434
rect 18732 44370 18788 44382
rect 18844 44996 18900 45006
rect 18844 44100 18900 44940
rect 18620 43540 18676 43550
rect 18508 43538 18676 43540
rect 18508 43486 18622 43538
rect 18674 43486 18676 43538
rect 18508 43484 18676 43486
rect 18620 43474 18676 43484
rect 18396 42130 18452 42140
rect 18732 42642 18788 42654
rect 18732 42590 18734 42642
rect 18786 42590 18788 42642
rect 18732 42084 18788 42590
rect 18732 42018 18788 42028
rect 18396 41972 18452 41982
rect 18396 41878 18452 41916
rect 18508 41186 18564 41198
rect 18508 41134 18510 41186
rect 18562 41134 18564 41186
rect 18284 40572 18452 40628
rect 18060 40404 18116 40414
rect 18284 40404 18340 40414
rect 18060 40310 18116 40348
rect 18172 40348 18284 40404
rect 17948 39788 18116 39844
rect 17836 39554 17892 39564
rect 17948 39618 18004 39630
rect 17948 39566 17950 39618
rect 18002 39566 18004 39618
rect 17948 38610 18004 39566
rect 17948 38558 17950 38610
rect 18002 38558 18004 38610
rect 17724 36036 17780 36204
rect 17388 35028 17444 35038
rect 17388 34914 17444 34972
rect 17388 34862 17390 34914
rect 17442 34862 17444 34914
rect 17388 34580 17444 34862
rect 17388 34514 17444 34524
rect 17276 32676 17332 33516
rect 17276 32610 17332 32620
rect 17388 33346 17444 33358
rect 17388 33294 17390 33346
rect 17442 33294 17444 33346
rect 17388 32788 17444 33294
rect 17388 32564 17444 32732
rect 17388 32498 17444 32508
rect 17276 31554 17332 31566
rect 17276 31502 17278 31554
rect 17330 31502 17332 31554
rect 17276 31220 17332 31502
rect 17500 31556 17556 35420
rect 17612 35980 17780 36036
rect 17836 38164 17892 38174
rect 17612 33572 17668 35980
rect 17724 35812 17780 35822
rect 17724 35718 17780 35756
rect 17724 33906 17780 33918
rect 17724 33854 17726 33906
rect 17778 33854 17780 33906
rect 17724 33796 17780 33854
rect 17724 33730 17780 33740
rect 17836 33906 17892 38108
rect 17948 38050 18004 38558
rect 18060 38164 18116 39788
rect 18060 38098 18116 38108
rect 17948 37998 17950 38050
rect 18002 37998 18004 38050
rect 17948 37986 18004 37998
rect 18060 37940 18116 37950
rect 18060 37490 18116 37884
rect 18060 37438 18062 37490
rect 18114 37438 18116 37490
rect 18060 37426 18116 37438
rect 18060 37044 18116 37054
rect 17948 36596 18004 36606
rect 17948 36502 18004 36540
rect 17948 36372 18004 36382
rect 17948 35812 18004 36316
rect 17948 35746 18004 35756
rect 17948 35476 18004 35486
rect 17948 35382 18004 35420
rect 18060 35140 18116 36988
rect 18172 36148 18228 40348
rect 18284 40310 18340 40348
rect 18284 39732 18340 39742
rect 18284 38834 18340 39676
rect 18284 38782 18286 38834
rect 18338 38782 18340 38834
rect 18284 38770 18340 38782
rect 18172 36082 18228 36092
rect 18284 38052 18340 38062
rect 18172 35812 18228 35822
rect 18172 35698 18228 35756
rect 18172 35646 18174 35698
rect 18226 35646 18228 35698
rect 18172 35634 18228 35646
rect 18060 35084 18228 35140
rect 17948 35028 18004 35038
rect 17948 35026 18116 35028
rect 17948 34974 17950 35026
rect 18002 34974 18116 35026
rect 17948 34972 18116 34974
rect 17948 34962 18004 34972
rect 18060 34356 18116 34972
rect 18060 34130 18116 34300
rect 18060 34078 18062 34130
rect 18114 34078 18116 34130
rect 18060 34066 18116 34078
rect 17836 33854 17838 33906
rect 17890 33854 17892 33906
rect 17612 33516 17780 33572
rect 17612 33124 17668 33134
rect 17612 33030 17668 33068
rect 17724 32900 17780 33516
rect 17500 31490 17556 31500
rect 17612 32844 17780 32900
rect 17276 31154 17332 31164
rect 17612 31108 17668 32844
rect 17724 32452 17780 32462
rect 17724 32004 17780 32396
rect 17724 31938 17780 31948
rect 17836 31892 17892 33854
rect 17836 31826 17892 31836
rect 18060 31892 18116 31902
rect 17836 31554 17892 31566
rect 17836 31502 17838 31554
rect 17890 31502 17892 31554
rect 17836 31332 17892 31502
rect 17836 31266 17892 31276
rect 17612 31052 17892 31108
rect 17836 30996 17892 31052
rect 17948 30996 18004 31006
rect 17836 30940 17948 30996
rect 17164 30436 17220 30940
rect 17948 30930 18004 30940
rect 17724 30884 17780 30894
rect 17724 30790 17780 30828
rect 17164 30370 17220 30380
rect 18060 30548 18116 31836
rect 18172 31668 18228 35084
rect 18284 35028 18340 37996
rect 18396 37828 18452 40572
rect 18508 40404 18564 41134
rect 18844 40516 18900 44044
rect 18956 43876 19012 48636
rect 19852 46788 19908 46798
rect 19852 46004 19908 46732
rect 19628 46002 19908 46004
rect 19628 45950 19854 46002
rect 19906 45950 19908 46002
rect 19628 45948 19908 45950
rect 18956 43762 19012 43820
rect 18956 43710 18958 43762
rect 19010 43710 19012 43762
rect 18956 43698 19012 43710
rect 19516 45332 19572 45342
rect 19516 45106 19572 45276
rect 19516 45054 19518 45106
rect 19570 45054 19572 45106
rect 19516 44324 19572 45054
rect 19628 45108 19684 45948
rect 19852 45938 19908 45948
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20188 45220 20244 49200
rect 22764 49028 22820 49038
rect 22204 46340 22260 46350
rect 22204 46002 22260 46284
rect 22204 45950 22206 46002
rect 22258 45950 22260 46002
rect 20636 45890 20692 45902
rect 20636 45838 20638 45890
rect 20690 45838 20692 45890
rect 20636 45332 20692 45838
rect 21532 45890 21588 45902
rect 21532 45838 21534 45890
rect 21586 45838 21588 45890
rect 20636 45266 20692 45276
rect 20860 45444 20916 45454
rect 20188 45154 20244 45164
rect 19628 45042 19684 45052
rect 19516 43708 19572 44268
rect 20300 44994 20356 45006
rect 20300 44942 20302 44994
rect 20354 44942 20356 44994
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 20188 43876 20244 43886
rect 19516 43652 19684 43708
rect 19628 43538 19684 43652
rect 19628 43486 19630 43538
rect 19682 43486 19684 43538
rect 19628 43474 19684 43486
rect 19404 43204 19460 43214
rect 18508 40338 18564 40348
rect 18620 40460 18900 40516
rect 18956 42756 19012 42766
rect 18956 42308 19012 42700
rect 18956 41186 19012 42252
rect 18956 41134 18958 41186
rect 19010 41134 19012 41186
rect 18396 37762 18452 37772
rect 18508 38276 18564 38286
rect 18396 37378 18452 37390
rect 18396 37326 18398 37378
rect 18450 37326 18452 37378
rect 18396 37268 18452 37326
rect 18396 37202 18452 37212
rect 18396 37044 18452 37054
rect 18396 35476 18452 36988
rect 18508 36260 18564 38220
rect 18620 37378 18676 40460
rect 18956 40404 19012 41134
rect 18844 40348 19012 40404
rect 18844 40290 18900 40348
rect 18844 40238 18846 40290
rect 18898 40238 18900 40290
rect 18844 40226 18900 40238
rect 18956 40292 19012 40348
rect 18956 40226 19012 40236
rect 19068 42084 19124 42094
rect 18732 39508 18788 39518
rect 18732 39414 18788 39452
rect 18844 39172 18900 39182
rect 18732 37938 18788 37950
rect 18732 37886 18734 37938
rect 18786 37886 18788 37938
rect 18732 37716 18788 37886
rect 18732 37650 18788 37660
rect 18620 37326 18622 37378
rect 18674 37326 18676 37378
rect 18620 37314 18676 37326
rect 18508 36204 18676 36260
rect 18508 36036 18564 36046
rect 18508 35812 18564 35980
rect 18508 35746 18564 35756
rect 18396 35382 18452 35420
rect 18284 34962 18340 34972
rect 18508 34804 18564 34814
rect 18284 34468 18340 34478
rect 18284 34130 18340 34412
rect 18284 34078 18286 34130
rect 18338 34078 18340 34130
rect 18284 34066 18340 34078
rect 18396 33906 18452 33918
rect 18396 33854 18398 33906
rect 18450 33854 18452 33906
rect 18396 33572 18452 33854
rect 18508 33908 18564 34748
rect 18508 33842 18564 33852
rect 18396 33506 18452 33516
rect 18620 33458 18676 36204
rect 18844 36148 18900 39116
rect 18956 37380 19012 37390
rect 18956 37266 19012 37324
rect 18956 37214 18958 37266
rect 19010 37214 19012 37266
rect 18956 36260 19012 37214
rect 18956 36194 19012 36204
rect 18620 33406 18622 33458
rect 18674 33406 18676 33458
rect 18620 33394 18676 33406
rect 18732 36092 18900 36148
rect 18732 33460 18788 36092
rect 18844 35924 18900 35934
rect 19068 35924 19124 42028
rect 19180 41858 19236 41870
rect 19180 41806 19182 41858
rect 19234 41806 19236 41858
rect 19180 41524 19236 41806
rect 19180 40402 19236 41468
rect 19180 40350 19182 40402
rect 19234 40350 19236 40402
rect 19180 40338 19236 40350
rect 19180 40180 19236 40190
rect 19180 39172 19236 40124
rect 19180 38834 19236 39116
rect 19180 38782 19182 38834
rect 19234 38782 19236 38834
rect 19180 38770 19236 38782
rect 19292 39844 19348 39854
rect 19292 38668 19348 39788
rect 18844 35922 19124 35924
rect 18844 35870 18846 35922
rect 18898 35870 19124 35922
rect 18844 35868 19124 35870
rect 19180 38612 19348 38668
rect 18844 35858 18900 35868
rect 19180 35476 19236 38612
rect 18732 33394 18788 33404
rect 18844 35420 19236 35476
rect 19292 36708 19348 36718
rect 19292 35698 19348 36652
rect 19292 35646 19294 35698
rect 19346 35646 19348 35698
rect 18284 33124 18340 33134
rect 18284 33122 18452 33124
rect 18284 33070 18286 33122
rect 18338 33070 18452 33122
rect 18284 33068 18452 33070
rect 18284 33058 18340 33068
rect 18284 32450 18340 32462
rect 18284 32398 18286 32450
rect 18338 32398 18340 32450
rect 18284 32004 18340 32398
rect 18284 31938 18340 31948
rect 18396 31892 18452 33068
rect 18508 33122 18564 33134
rect 18508 33070 18510 33122
rect 18562 33070 18564 33122
rect 18508 32564 18564 33070
rect 18732 33124 18788 33134
rect 18732 33030 18788 33068
rect 18844 32786 18900 35420
rect 19292 35364 19348 35646
rect 19180 35308 19348 35364
rect 19180 34130 19236 35308
rect 19404 34244 19460 43148
rect 20188 42868 20244 43820
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19516 41972 19572 41982
rect 19516 37492 19572 41916
rect 19964 41860 20020 41870
rect 19964 41188 20020 41804
rect 19964 41056 20020 41132
rect 19628 40852 19684 40862
rect 19628 40626 19684 40796
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19628 40574 19630 40626
rect 19682 40574 19684 40626
rect 19628 40562 19684 40574
rect 19964 40402 20020 40414
rect 19964 40350 19966 40402
rect 20018 40350 20020 40402
rect 19964 39396 20020 40350
rect 19628 39340 20020 39396
rect 19628 39060 19684 39340
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19628 39004 19908 39060
rect 19740 38836 19796 38846
rect 19628 38834 19796 38836
rect 19628 38782 19742 38834
rect 19794 38782 19796 38834
rect 19628 38780 19796 38782
rect 19628 38052 19684 38780
rect 19740 38770 19796 38780
rect 19628 37986 19684 37996
rect 19852 38724 19908 39004
rect 19852 37828 19908 38668
rect 19516 37154 19572 37436
rect 19516 37102 19518 37154
rect 19570 37102 19572 37154
rect 19516 37090 19572 37102
rect 19628 37772 19908 37828
rect 19404 34178 19460 34188
rect 19516 36484 19572 36494
rect 19180 34078 19182 34130
rect 19234 34078 19236 34130
rect 19180 34066 19236 34078
rect 19292 34132 19348 34142
rect 18844 32734 18846 32786
rect 18898 32734 18900 32786
rect 18844 32722 18900 32734
rect 19292 32676 19348 34076
rect 19404 33684 19460 33694
rect 19404 33570 19460 33628
rect 19404 33518 19406 33570
rect 19458 33518 19460 33570
rect 19404 33506 19460 33518
rect 19404 32676 19460 32686
rect 19292 32674 19460 32676
rect 19292 32622 19406 32674
rect 19458 32622 19460 32674
rect 19292 32620 19460 32622
rect 19404 32610 19460 32620
rect 19516 32564 19572 36428
rect 19628 32788 19684 37772
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 20076 36484 20132 36494
rect 20076 36390 20132 36428
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 20076 35812 20132 35822
rect 20076 35718 20132 35756
rect 20076 34804 20132 34814
rect 20076 34710 20132 34748
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19852 34244 19908 34254
rect 19852 34018 19908 34188
rect 19852 33966 19854 34018
rect 19906 33966 19908 34018
rect 19852 33572 19908 33966
rect 19852 33506 19908 33516
rect 19740 33460 19796 33470
rect 19740 33346 19796 33404
rect 20076 33460 20132 33470
rect 20076 33366 20132 33404
rect 19740 33294 19742 33346
rect 19794 33294 19796 33346
rect 19740 33282 19796 33294
rect 20188 33236 20244 42812
rect 20300 39956 20356 44942
rect 20412 44548 20468 44558
rect 20412 43426 20468 44492
rect 20860 44434 20916 45388
rect 21532 45332 21588 45838
rect 20860 44382 20862 44434
rect 20914 44382 20916 44434
rect 20860 44370 20916 44382
rect 21196 44660 21252 44670
rect 21196 43708 21252 44604
rect 21532 44324 21588 45276
rect 21868 44884 21924 44894
rect 21644 44324 21700 44334
rect 21532 44322 21700 44324
rect 21532 44270 21646 44322
rect 21698 44270 21700 44322
rect 21532 44268 21700 44270
rect 21644 44258 21700 44268
rect 21196 43652 21364 43708
rect 20412 43374 20414 43426
rect 20466 43374 20468 43426
rect 20412 42868 20468 43374
rect 20412 42802 20468 42812
rect 20860 42868 20916 42878
rect 20860 42774 20916 42812
rect 21196 42308 21252 42318
rect 20972 41412 21028 41422
rect 20860 41076 20916 41086
rect 20860 40982 20916 41020
rect 20748 40964 20804 40974
rect 20636 40962 20804 40964
rect 20636 40910 20750 40962
rect 20802 40910 20804 40962
rect 20636 40908 20804 40910
rect 20412 40516 20468 40526
rect 20412 40180 20468 40460
rect 20412 40114 20468 40124
rect 20524 40292 20580 40302
rect 20300 39890 20356 39900
rect 20188 33170 20244 33180
rect 20412 38946 20468 38958
rect 20412 38894 20414 38946
rect 20466 38894 20468 38946
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19628 32732 20132 32788
rect 19740 32564 19796 32574
rect 18508 32508 18788 32564
rect 19516 32562 19796 32564
rect 19516 32510 19742 32562
rect 19794 32510 19796 32562
rect 19516 32508 19796 32510
rect 18508 32340 18564 32350
rect 18508 32246 18564 32284
rect 18396 31826 18452 31836
rect 18620 31892 18676 31902
rect 18508 31780 18564 31790
rect 18508 31686 18564 31724
rect 18284 31668 18340 31678
rect 18172 31666 18340 31668
rect 18172 31614 18286 31666
rect 18338 31614 18340 31666
rect 18172 31612 18340 31614
rect 18284 31602 18340 31612
rect 18508 31556 18564 31566
rect 18508 31218 18564 31500
rect 18508 31166 18510 31218
rect 18562 31166 18564 31218
rect 18508 31154 18564 31166
rect 18172 30996 18228 31006
rect 18172 30902 18228 30940
rect 17276 30324 17332 30334
rect 17276 30230 17332 30268
rect 17836 30324 17892 30334
rect 17836 30230 17892 30268
rect 18060 26908 18116 30492
rect 18284 30212 18340 30222
rect 18620 30212 18676 31836
rect 18732 31668 18788 32508
rect 19516 32338 19572 32350
rect 19516 32286 19518 32338
rect 19570 32286 19572 32338
rect 19516 32116 19572 32286
rect 19516 32050 19572 32060
rect 19180 31892 19236 31902
rect 19180 31778 19236 31836
rect 19180 31726 19182 31778
rect 19234 31726 19236 31778
rect 19180 31714 19236 31726
rect 18732 31602 18788 31612
rect 19068 31668 19124 31678
rect 19068 31332 19124 31612
rect 19740 31668 19796 32508
rect 19964 32338 20020 32350
rect 19964 32286 19966 32338
rect 20018 32286 20020 32338
rect 19964 32004 20020 32286
rect 19964 31938 20020 31948
rect 20076 31780 20132 32732
rect 20188 32562 20244 32574
rect 20188 32510 20190 32562
rect 20242 32510 20244 32562
rect 20188 32004 20244 32510
rect 20412 32116 20468 38894
rect 20524 38834 20580 40236
rect 20636 39396 20692 40908
rect 20748 40898 20804 40908
rect 20748 40404 20804 40414
rect 20748 40310 20804 40348
rect 20860 39732 20916 39742
rect 20860 39638 20916 39676
rect 20636 39330 20692 39340
rect 20524 38782 20526 38834
rect 20578 38782 20580 38834
rect 20524 36484 20580 38782
rect 20972 38836 21028 41356
rect 21196 41188 21252 42252
rect 21196 40628 21252 41132
rect 21196 40402 21252 40572
rect 21196 40350 21198 40402
rect 21250 40350 21252 40402
rect 21196 40338 21252 40350
rect 21196 39956 21252 39966
rect 21196 39396 21252 39900
rect 21196 39330 21252 39340
rect 21084 38836 21140 38846
rect 20972 38834 21140 38836
rect 20972 38782 21086 38834
rect 21138 38782 21140 38834
rect 20972 38780 21140 38782
rect 21084 38668 21140 38780
rect 21084 38612 21252 38668
rect 20860 38164 20916 38174
rect 20860 38070 20916 38108
rect 20524 36418 20580 36428
rect 20748 38052 20804 38062
rect 20748 36708 20804 37996
rect 20748 36482 20804 36652
rect 20748 36430 20750 36482
rect 20802 36430 20804 36482
rect 20748 34914 20804 36430
rect 20748 34862 20750 34914
rect 20802 34862 20804 34914
rect 20748 34850 20804 34862
rect 21084 35700 21140 35710
rect 20860 33572 20916 33582
rect 20860 33458 20916 33516
rect 20860 33406 20862 33458
rect 20914 33406 20916 33458
rect 20860 33394 20916 33406
rect 20412 32050 20468 32060
rect 20636 33236 20692 33246
rect 20188 31938 20244 31948
rect 20300 31836 20580 31892
rect 20188 31780 20244 31790
rect 20076 31778 20244 31780
rect 20076 31726 20190 31778
rect 20242 31726 20244 31778
rect 20076 31724 20244 31726
rect 19740 31602 19796 31612
rect 19068 31266 19124 31276
rect 19404 31556 19460 31566
rect 19068 31108 19124 31118
rect 19404 31108 19460 31500
rect 19516 31556 19572 31566
rect 19516 31554 19684 31556
rect 19516 31502 19518 31554
rect 19570 31502 19684 31554
rect 19516 31500 19684 31502
rect 19516 31490 19572 31500
rect 19516 31108 19572 31118
rect 19068 30772 19124 31052
rect 19068 30706 19124 30716
rect 19292 31106 19572 31108
rect 19292 31054 19518 31106
rect 19570 31054 19572 31106
rect 19292 31052 19572 31054
rect 18284 30210 18676 30212
rect 18284 30158 18286 30210
rect 18338 30158 18676 30210
rect 18284 30156 18676 30158
rect 18284 30146 18340 30156
rect 18620 29652 18676 30156
rect 19068 30548 19124 30558
rect 18732 29986 18788 29998
rect 18732 29934 18734 29986
rect 18786 29934 18788 29986
rect 18732 29876 18788 29934
rect 18732 29810 18788 29820
rect 19068 29652 19124 30492
rect 19180 30212 19236 30222
rect 19180 30118 19236 30156
rect 19180 29652 19236 29662
rect 19068 29650 19236 29652
rect 19068 29598 19182 29650
rect 19234 29598 19236 29650
rect 19068 29596 19236 29598
rect 18620 29586 18676 29596
rect 19180 29586 19236 29596
rect 19292 26908 19348 31052
rect 19516 31042 19572 31052
rect 19628 30548 19684 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19740 31220 19796 31230
rect 19740 31126 19796 31164
rect 19628 30482 19684 30492
rect 19740 30772 19796 30782
rect 19628 30324 19684 30334
rect 19740 30324 19796 30716
rect 19628 30322 19796 30324
rect 19628 30270 19630 30322
rect 19682 30270 19796 30322
rect 19628 30268 19796 30270
rect 19852 30770 19908 30782
rect 19852 30718 19854 30770
rect 19906 30718 19908 30770
rect 19628 30258 19684 30268
rect 19852 30100 19908 30718
rect 20188 30324 20244 31724
rect 20300 31778 20356 31836
rect 20300 31726 20302 31778
rect 20354 31726 20356 31778
rect 20300 31714 20356 31726
rect 20412 31666 20468 31678
rect 20412 31614 20414 31666
rect 20466 31614 20468 31666
rect 20412 30996 20468 31614
rect 20076 30268 20244 30324
rect 20300 30940 20468 30996
rect 20524 30996 20580 31836
rect 20076 30210 20132 30268
rect 20076 30158 20078 30210
rect 20130 30158 20132 30210
rect 20076 30146 20132 30158
rect 19852 30034 19908 30044
rect 20300 29988 20356 30940
rect 20524 30930 20580 30940
rect 20300 29922 20356 29932
rect 20412 30770 20468 30782
rect 20412 30718 20414 30770
rect 20466 30718 20468 30770
rect 20412 30660 20468 30718
rect 20524 30772 20580 30782
rect 20524 30678 20580 30716
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 18060 26852 18452 26908
rect 16716 26338 16772 26348
rect 18396 24724 18452 26852
rect 18396 24658 18452 24668
rect 19068 26852 19348 26908
rect 19404 29652 19460 29662
rect 19068 24052 19124 26852
rect 19068 23986 19124 23996
rect 16156 16706 16212 16716
rect 15036 16370 15092 16380
rect 6636 15026 6692 15036
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 1820 14306 1876 14318
rect 1820 14254 1822 14306
rect 1874 14254 1876 14306
rect 1820 14196 1876 14254
rect 1820 14130 1876 14140
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 19404 11508 19460 29596
rect 19740 29652 19796 29662
rect 19740 29558 19796 29596
rect 20300 29314 20356 29326
rect 20300 29262 20302 29314
rect 20354 29262 20356 29314
rect 20300 29202 20356 29262
rect 20300 29150 20302 29202
rect 20354 29150 20356 29202
rect 20300 29138 20356 29150
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20412 27412 20468 30604
rect 20524 29986 20580 29998
rect 20524 29934 20526 29986
rect 20578 29934 20580 29986
rect 20524 29876 20580 29934
rect 20524 29810 20580 29820
rect 20636 29202 20692 33180
rect 20860 33124 20916 33134
rect 20748 32338 20804 32350
rect 20748 32286 20750 32338
rect 20802 32286 20804 32338
rect 20748 32228 20804 32286
rect 20748 32004 20804 32172
rect 20748 31938 20804 31948
rect 20860 31554 20916 33068
rect 21084 32674 21140 35644
rect 21084 32622 21086 32674
rect 21138 32622 21140 32674
rect 21084 32610 21140 32622
rect 20860 31502 20862 31554
rect 20914 31502 20916 31554
rect 20860 31332 20916 31502
rect 20972 32562 21028 32574
rect 20972 32510 20974 32562
rect 21026 32510 21028 32562
rect 20972 32228 21028 32510
rect 20972 31556 21028 32172
rect 20972 31490 21028 31500
rect 21084 32116 21140 32126
rect 20860 31276 21028 31332
rect 20748 30770 20804 30782
rect 20748 30718 20750 30770
rect 20802 30718 20804 30770
rect 20748 30548 20804 30718
rect 20748 30482 20804 30492
rect 20860 30770 20916 30782
rect 20860 30718 20862 30770
rect 20914 30718 20916 30770
rect 20860 30436 20916 30718
rect 20860 30370 20916 30380
rect 20748 30324 20804 30334
rect 20748 29650 20804 30268
rect 20860 30212 20916 30222
rect 20860 30098 20916 30156
rect 20860 30046 20862 30098
rect 20914 30046 20916 30098
rect 20860 29876 20916 30046
rect 20860 29810 20916 29820
rect 20972 29764 21028 31276
rect 20972 29698 21028 29708
rect 20748 29598 20750 29650
rect 20802 29598 20804 29650
rect 20748 29586 20804 29598
rect 20860 29652 20916 29662
rect 20860 29316 20916 29596
rect 21084 29540 21140 32060
rect 21196 30996 21252 38612
rect 21308 33572 21364 43652
rect 21644 42866 21700 42878
rect 21644 42814 21646 42866
rect 21698 42814 21700 42866
rect 21644 42756 21700 42814
rect 21644 42690 21700 42700
rect 21420 41858 21476 41870
rect 21420 41806 21422 41858
rect 21474 41806 21476 41858
rect 21420 41748 21476 41806
rect 21420 41682 21476 41692
rect 21756 41188 21812 41198
rect 21868 41188 21924 44828
rect 22204 44436 22260 45950
rect 22428 44996 22484 45006
rect 22428 44994 22596 44996
rect 22428 44942 22430 44994
rect 22482 44942 22596 44994
rect 22428 44940 22596 44942
rect 22428 44930 22484 44940
rect 22204 44370 22260 44380
rect 22428 44772 22484 44782
rect 22428 44434 22484 44716
rect 22428 44382 22430 44434
rect 22482 44382 22484 44434
rect 22428 44370 22484 44382
rect 22540 43988 22596 44940
rect 22540 43708 22596 43932
rect 22204 43652 22260 43662
rect 21756 41186 21924 41188
rect 21756 41134 21758 41186
rect 21810 41134 21924 41186
rect 21756 41132 21924 41134
rect 21980 43092 22036 43102
rect 21756 41122 21812 41132
rect 21420 40628 21476 40638
rect 21420 38946 21476 40572
rect 21420 38894 21422 38946
rect 21474 38894 21476 38946
rect 21420 38882 21476 38894
rect 21532 40404 21588 40414
rect 21532 38668 21588 40348
rect 21420 38612 21588 38668
rect 21644 39618 21700 39630
rect 21644 39566 21646 39618
rect 21698 39566 21700 39618
rect 21644 38612 21700 39566
rect 21980 39060 22036 43036
rect 22092 41972 22148 42010
rect 22092 41906 22148 41916
rect 22092 41748 22148 41758
rect 22204 41748 22260 43596
rect 22428 43652 22596 43708
rect 22652 44884 22708 44894
rect 22652 43652 22708 44828
rect 22148 41692 22260 41748
rect 22316 41972 22372 41982
rect 22092 40180 22148 41692
rect 22204 40516 22260 40526
rect 22204 40402 22260 40460
rect 22204 40350 22206 40402
rect 22258 40350 22260 40402
rect 22204 40338 22260 40350
rect 22092 40124 22260 40180
rect 21420 36484 21476 38612
rect 21644 38052 21700 38556
rect 21644 37958 21700 37996
rect 21868 39004 22036 39060
rect 21868 37940 21924 39004
rect 21980 38834 22036 38846
rect 21980 38782 21982 38834
rect 22034 38782 22036 38834
rect 21980 38612 22036 38782
rect 21980 38546 22036 38556
rect 21644 37156 21700 37166
rect 21644 37154 21812 37156
rect 21644 37102 21646 37154
rect 21698 37102 21812 37154
rect 21644 37100 21812 37102
rect 21644 37090 21700 37100
rect 21644 36596 21700 36606
rect 21644 36502 21700 36540
rect 21420 36428 21588 36484
rect 21308 32788 21364 33516
rect 21308 32722 21364 32732
rect 21532 32564 21588 36428
rect 21756 35140 21812 37100
rect 21756 35074 21812 35084
rect 21644 35028 21700 35038
rect 21644 34934 21700 34972
rect 21868 33684 21924 37884
rect 22092 37828 22148 37838
rect 21980 37716 22036 37726
rect 21980 36820 22036 37660
rect 21980 36754 22036 36764
rect 21980 35140 22036 35150
rect 21980 34018 22036 35084
rect 21980 33966 21982 34018
rect 22034 33966 22036 34018
rect 21980 33796 22036 33966
rect 21980 33730 22036 33740
rect 21756 33628 21924 33684
rect 21756 33012 21812 33628
rect 21868 33458 21924 33470
rect 21868 33406 21870 33458
rect 21922 33406 21924 33458
rect 21868 33236 21924 33406
rect 21868 33170 21924 33180
rect 21980 33346 22036 33358
rect 21980 33294 21982 33346
rect 22034 33294 22036 33346
rect 21756 32956 21924 33012
rect 21532 32508 21700 32564
rect 21196 30930 21252 30940
rect 21308 32452 21364 32462
rect 21308 32338 21364 32396
rect 21308 32286 21310 32338
rect 21362 32286 21364 32338
rect 21308 30100 21364 32286
rect 21532 32340 21588 32350
rect 21532 32246 21588 32284
rect 21644 32116 21700 32508
rect 21532 32060 21700 32116
rect 21532 31444 21588 32060
rect 21532 31378 21588 31388
rect 21644 31892 21700 31902
rect 21644 31778 21700 31836
rect 21644 31726 21646 31778
rect 21698 31726 21700 31778
rect 21308 30034 21364 30044
rect 21532 30770 21588 30782
rect 21532 30718 21534 30770
rect 21586 30718 21588 30770
rect 21196 29876 21252 29886
rect 21196 29650 21252 29820
rect 21196 29598 21198 29650
rect 21250 29598 21252 29650
rect 21196 29586 21252 29598
rect 21084 29474 21140 29484
rect 20860 29250 20916 29260
rect 20636 29150 20638 29202
rect 20690 29150 20692 29202
rect 20636 29138 20692 29150
rect 21532 27860 21588 30718
rect 21644 30772 21700 31726
rect 21868 31890 21924 32956
rect 21980 32564 22036 33294
rect 21980 32498 22036 32508
rect 21868 31838 21870 31890
rect 21922 31838 21924 31890
rect 21868 31220 21924 31838
rect 22092 31892 22148 37772
rect 22204 37604 22260 40124
rect 22204 35586 22260 37548
rect 22316 38612 22372 41916
rect 22428 41636 22484 43652
rect 22652 43586 22708 43596
rect 22540 43428 22596 43438
rect 22540 43426 22708 43428
rect 22540 43374 22542 43426
rect 22594 43374 22708 43426
rect 22540 43372 22708 43374
rect 22540 43362 22596 43372
rect 22652 43204 22708 43372
rect 22652 43138 22708 43148
rect 22764 42082 22820 48972
rect 22988 48804 23044 48814
rect 22988 48710 23044 48748
rect 22764 42030 22766 42082
rect 22818 42030 22820 42082
rect 22428 41580 22596 41636
rect 22316 37266 22372 38556
rect 22428 39506 22484 39518
rect 22428 39454 22430 39506
rect 22482 39454 22484 39506
rect 22428 38164 22484 39454
rect 22540 38724 22596 41580
rect 22652 41186 22708 41198
rect 22652 41134 22654 41186
rect 22706 41134 22708 41186
rect 22652 40292 22708 41134
rect 22652 40226 22708 40236
rect 22764 40068 22820 42030
rect 22876 46004 22932 46014
rect 22876 42084 22932 45948
rect 22988 45220 23044 45230
rect 22988 45126 23044 45164
rect 22876 41524 22932 42028
rect 23100 45106 23156 45118
rect 23100 45054 23102 45106
rect 23154 45054 23156 45106
rect 23100 42084 23156 45054
rect 23100 42018 23156 42028
rect 23212 41858 23268 49308
rect 23520 49200 23632 49800
rect 24892 49700 24948 49710
rect 23660 47794 23716 47806
rect 23660 47742 23662 47794
rect 23714 47742 23716 47794
rect 23212 41806 23214 41858
rect 23266 41806 23268 41858
rect 22876 41468 23044 41524
rect 22988 40514 23044 41468
rect 22988 40462 22990 40514
rect 23042 40462 23044 40514
rect 22988 40450 23044 40462
rect 22764 40002 22820 40012
rect 22876 40402 22932 40414
rect 22876 40350 22878 40402
rect 22930 40350 22932 40402
rect 22764 38724 22820 38734
rect 22540 38722 22820 38724
rect 22540 38670 22766 38722
rect 22818 38670 22820 38722
rect 22540 38668 22820 38670
rect 22428 38098 22484 38108
rect 22316 37214 22318 37266
rect 22370 37214 22372 37266
rect 22316 37156 22372 37214
rect 22316 37090 22372 37100
rect 22428 37940 22484 37950
rect 22428 37044 22484 37884
rect 22764 37716 22820 38668
rect 22764 37650 22820 37660
rect 22428 36978 22484 36988
rect 22540 37380 22596 37390
rect 22204 35534 22206 35586
rect 22258 35534 22260 35586
rect 22204 35522 22260 35534
rect 22428 35028 22484 35038
rect 22204 33572 22260 33582
rect 22204 32786 22260 33516
rect 22204 32734 22206 32786
rect 22258 32734 22260 32786
rect 22204 32722 22260 32734
rect 22316 33460 22372 33470
rect 22316 32786 22372 33404
rect 22428 33124 22484 34972
rect 22540 33348 22596 37324
rect 22876 37268 22932 40350
rect 22652 37212 22932 37268
rect 22988 40292 23044 40302
rect 22652 33684 22708 37212
rect 22988 37044 23044 40236
rect 22876 36988 23044 37044
rect 23100 37044 23156 37054
rect 22876 35922 22932 36988
rect 23100 36950 23156 36988
rect 22876 35870 22878 35922
rect 22930 35870 22932 35922
rect 22876 35858 22932 35870
rect 23212 35812 23268 41806
rect 23324 47460 23380 47470
rect 23324 43538 23380 47404
rect 23660 47348 23716 47742
rect 23996 47794 24052 47806
rect 23996 47742 23998 47794
rect 24050 47742 24052 47794
rect 23660 47282 23716 47292
rect 23884 47348 23940 47358
rect 23772 45106 23828 45118
rect 23772 45054 23774 45106
rect 23826 45054 23828 45106
rect 23324 43486 23326 43538
rect 23378 43486 23380 43538
rect 23324 41860 23380 43486
rect 23660 44100 23716 44110
rect 23548 43428 23604 43438
rect 23548 43314 23604 43372
rect 23660 43426 23716 44044
rect 23660 43374 23662 43426
rect 23714 43374 23716 43426
rect 23660 43362 23716 43374
rect 23548 43262 23550 43314
rect 23602 43262 23604 43314
rect 23548 42756 23604 43262
rect 23772 43092 23828 45054
rect 23772 43026 23828 43036
rect 23772 42868 23828 42878
rect 23884 42868 23940 47292
rect 23772 42866 23940 42868
rect 23772 42814 23774 42866
rect 23826 42814 23940 42866
rect 23772 42812 23940 42814
rect 23772 42802 23828 42812
rect 23548 42700 23716 42756
rect 23324 41794 23380 41804
rect 23548 42532 23604 42542
rect 23436 40740 23492 40750
rect 23100 35756 23268 35812
rect 23324 38052 23380 38062
rect 22876 35698 22932 35710
rect 22876 35646 22878 35698
rect 22930 35646 22932 35698
rect 22876 33908 22932 35646
rect 23100 35364 23156 35756
rect 23324 35698 23380 37996
rect 23324 35646 23326 35698
rect 23378 35646 23380 35698
rect 23324 35634 23380 35646
rect 23436 37828 23492 40684
rect 23548 40626 23604 42476
rect 23660 41972 23716 42700
rect 23884 42084 23940 42094
rect 23660 41916 23828 41972
rect 23660 41298 23716 41310
rect 23660 41246 23662 41298
rect 23714 41246 23716 41298
rect 23660 41188 23716 41246
rect 23660 41122 23716 41132
rect 23548 40574 23550 40626
rect 23602 40574 23604 40626
rect 23548 40562 23604 40574
rect 23772 38668 23828 41916
rect 23436 35476 23492 37772
rect 23324 35420 23492 35476
rect 23660 38612 23828 38668
rect 23100 35308 23268 35364
rect 23100 34132 23156 34142
rect 23100 34038 23156 34076
rect 22876 33842 22932 33852
rect 22988 33796 23044 33806
rect 22988 33684 23044 33740
rect 22652 33628 22820 33684
rect 22652 33348 22708 33358
rect 22540 33346 22708 33348
rect 22540 33294 22654 33346
rect 22706 33294 22708 33346
rect 22540 33292 22708 33294
rect 22652 33282 22708 33292
rect 22428 33068 22708 33124
rect 22316 32734 22318 32786
rect 22370 32734 22372 32786
rect 22316 32722 22372 32734
rect 22428 32674 22484 32686
rect 22428 32622 22430 32674
rect 22482 32622 22484 32674
rect 22092 31836 22372 31892
rect 22204 31556 22260 31566
rect 22204 31462 22260 31500
rect 22316 31444 22372 31836
rect 22428 31668 22484 32622
rect 22540 32676 22596 32686
rect 22540 32582 22596 32620
rect 22652 32004 22708 33068
rect 22652 31938 22708 31948
rect 22764 31892 22820 33628
rect 22876 33628 23044 33684
rect 22876 32676 22932 33628
rect 23212 33460 23268 35308
rect 23212 33394 23268 33404
rect 23324 33348 23380 35420
rect 23548 35252 23604 35262
rect 23548 34804 23604 35196
rect 23548 34738 23604 34748
rect 23436 34018 23492 34030
rect 23436 33966 23438 34018
rect 23490 33966 23492 34018
rect 23436 33796 23492 33966
rect 23548 33908 23604 33918
rect 23548 33814 23604 33852
rect 23436 33730 23492 33740
rect 23660 33796 23716 38612
rect 23884 37828 23940 42028
rect 23772 37772 23940 37828
rect 23772 37156 23828 37772
rect 23884 37604 23940 37614
rect 23884 37378 23940 37548
rect 23884 37326 23886 37378
rect 23938 37326 23940 37378
rect 23884 37314 23940 37326
rect 23772 37100 23940 37156
rect 23772 36596 23828 36606
rect 23772 36502 23828 36540
rect 23884 35700 23940 37100
rect 23996 37154 24052 47742
rect 24220 47124 24276 47134
rect 24108 43540 24164 43550
rect 24108 43446 24164 43484
rect 24108 41970 24164 41982
rect 24108 41918 24110 41970
rect 24162 41918 24164 41970
rect 24108 38052 24164 41918
rect 24220 41972 24276 47068
rect 24332 46002 24388 46014
rect 24332 45950 24334 46002
rect 24386 45950 24388 46002
rect 24332 42196 24388 45950
rect 24892 45220 24948 49644
rect 25536 49200 25648 49800
rect 25844 49756 25956 49812
rect 25788 49746 25844 49756
rect 25788 49476 25844 49486
rect 25564 49028 25620 49038
rect 25564 48934 25620 48972
rect 25788 49028 25844 49420
rect 25788 46002 25844 48972
rect 25788 45950 25790 46002
rect 25842 45950 25844 46002
rect 25788 45938 25844 45950
rect 24444 45106 24500 45118
rect 24444 45054 24446 45106
rect 24498 45054 24500 45106
rect 24444 43428 24500 45054
rect 24892 44996 24948 45164
rect 25676 45780 25732 45790
rect 24892 44994 25060 44996
rect 24892 44942 24894 44994
rect 24946 44942 25060 44994
rect 24892 44940 25060 44942
rect 24892 44930 24948 44940
rect 24556 44884 24612 44894
rect 24556 44882 24724 44884
rect 24556 44830 24558 44882
rect 24610 44830 24724 44882
rect 24556 44828 24724 44830
rect 24556 44818 24612 44828
rect 24556 44436 24612 44446
rect 24556 44342 24612 44380
rect 24556 43540 24612 43550
rect 24556 43446 24612 43484
rect 24444 43362 24500 43372
rect 24556 42756 24612 42766
rect 24556 42662 24612 42700
rect 24332 42140 24612 42196
rect 24332 41972 24388 41982
rect 24220 41970 24388 41972
rect 24220 41918 24334 41970
rect 24386 41918 24388 41970
rect 24220 41916 24388 41918
rect 24220 41300 24276 41310
rect 24220 41186 24276 41244
rect 24220 41134 24222 41186
rect 24274 41134 24276 41186
rect 24220 41122 24276 41134
rect 24332 39844 24388 41916
rect 24444 41972 24500 41982
rect 24444 41746 24500 41916
rect 24444 41694 24446 41746
rect 24498 41694 24500 41746
rect 24444 41682 24500 41694
rect 24556 40964 24612 42140
rect 24668 41186 24724 44828
rect 24780 44772 24836 44782
rect 24780 43708 24836 44716
rect 25004 44772 25060 44940
rect 25004 44706 25060 44716
rect 25340 44436 25396 44446
rect 25228 44322 25284 44334
rect 25228 44270 25230 44322
rect 25282 44270 25284 44322
rect 25228 43708 25284 44270
rect 24780 43652 24948 43708
rect 24668 41134 24670 41186
rect 24722 41134 24724 41186
rect 24668 41122 24724 41134
rect 24556 40908 24724 40964
rect 24556 40740 24612 40750
rect 24444 40514 24500 40526
rect 24444 40462 24446 40514
rect 24498 40462 24500 40514
rect 24444 40404 24500 40462
rect 24444 40338 24500 40348
rect 24556 40402 24612 40684
rect 24556 40350 24558 40402
rect 24610 40350 24612 40402
rect 24556 40338 24612 40350
rect 24108 37986 24164 37996
rect 24220 39788 24388 39844
rect 23996 37102 23998 37154
rect 24050 37102 24052 37154
rect 23996 37090 24052 37102
rect 24220 36932 24276 39788
rect 24556 39730 24612 39742
rect 24556 39678 24558 39730
rect 24610 39678 24612 39730
rect 24556 39620 24612 39678
rect 24444 39508 24500 39518
rect 24444 38948 24500 39452
rect 24556 39172 24612 39564
rect 24556 39106 24612 39116
rect 24668 38948 24724 40908
rect 24892 39508 24948 43652
rect 25116 43652 25284 43708
rect 25116 42866 25172 43652
rect 25116 42814 25118 42866
rect 25170 42814 25172 42866
rect 25116 42756 25172 42814
rect 25116 42196 25172 42700
rect 25340 42980 25396 44380
rect 25676 43426 25732 45724
rect 25676 43374 25678 43426
rect 25730 43374 25732 43426
rect 25676 43362 25732 43374
rect 25788 45106 25844 45118
rect 25788 45054 25790 45106
rect 25842 45054 25844 45106
rect 25116 42130 25172 42140
rect 25228 42532 25284 42542
rect 25116 40404 25172 40414
rect 25116 39732 25172 40348
rect 25228 39956 25284 42476
rect 25340 41300 25396 42924
rect 25788 42420 25844 45054
rect 25900 44436 25956 49756
rect 26012 49588 26068 49598
rect 26124 49588 26180 49756
rect 26068 49532 26180 49588
rect 26236 49588 26292 49598
rect 26012 49522 26068 49532
rect 26012 49140 26068 49150
rect 26236 49140 26292 49532
rect 26068 49084 26292 49140
rect 26572 49252 26628 49262
rect 26880 49200 26992 49800
rect 28896 49200 29008 49800
rect 30912 49200 31024 49800
rect 31948 49252 32004 49262
rect 26012 49074 26068 49084
rect 26460 49028 26516 49038
rect 26460 48934 26516 48972
rect 26012 48804 26068 48814
rect 26012 45892 26068 48748
rect 26572 48020 26628 49196
rect 26348 46002 26404 46014
rect 26348 45950 26350 46002
rect 26402 45950 26404 46002
rect 26012 45890 26180 45892
rect 26012 45838 26014 45890
rect 26066 45838 26180 45890
rect 26012 45836 26180 45838
rect 26012 45826 26068 45836
rect 25900 44304 25956 44380
rect 26012 45218 26068 45230
rect 26012 45166 26014 45218
rect 26066 45166 26068 45218
rect 25788 42354 25844 42364
rect 25788 42196 25844 42206
rect 25788 41970 25844 42140
rect 25788 41918 25790 41970
rect 25842 41918 25844 41970
rect 25788 41906 25844 41918
rect 25340 41298 25508 41300
rect 25340 41246 25342 41298
rect 25394 41246 25508 41298
rect 25340 41244 25508 41246
rect 25340 41234 25396 41244
rect 25228 39890 25284 39900
rect 25340 40180 25396 40190
rect 24892 39442 24948 39452
rect 25004 39730 25172 39732
rect 25004 39678 25118 39730
rect 25170 39678 25172 39730
rect 25004 39676 25172 39678
rect 24444 38892 24612 38948
rect 24444 38724 24500 38734
rect 24220 36866 24276 36876
rect 24332 38612 24500 38668
rect 24332 36036 24388 38612
rect 24556 38162 24612 38892
rect 24668 38882 24724 38892
rect 24892 38724 24948 38734
rect 24892 38630 24948 38668
rect 24556 38110 24558 38162
rect 24610 38110 24612 38162
rect 24108 35980 24388 36036
rect 24444 37156 24500 37166
rect 24444 36482 24500 37100
rect 24556 36708 24612 38110
rect 25004 37940 25060 39676
rect 25116 39666 25172 39676
rect 25004 37874 25060 37884
rect 25228 38052 25284 38062
rect 25340 38052 25396 40124
rect 25228 38050 25396 38052
rect 25228 37998 25230 38050
rect 25282 37998 25396 38050
rect 25228 37996 25396 37998
rect 25116 37604 25172 37614
rect 24556 36642 24612 36652
rect 24668 37044 24724 37054
rect 24444 36430 24446 36482
rect 24498 36430 24500 36482
rect 23996 35700 24052 35710
rect 23884 35698 24052 35700
rect 23884 35646 23998 35698
rect 24050 35646 24052 35698
rect 23884 35644 24052 35646
rect 23884 35028 23940 35644
rect 23996 35634 24052 35644
rect 23772 34804 23828 34814
rect 23772 34710 23828 34748
rect 23884 34580 23940 34972
rect 23884 34514 23940 34524
rect 23996 35364 24052 35374
rect 23660 33730 23716 33740
rect 23772 33572 23828 33582
rect 23772 33478 23828 33516
rect 23660 33460 23716 33470
rect 23324 33346 23492 33348
rect 23324 33294 23326 33346
rect 23378 33294 23492 33346
rect 23324 33292 23492 33294
rect 23324 33282 23380 33292
rect 23212 33236 23268 33246
rect 22876 32610 22932 32620
rect 23100 33234 23268 33236
rect 23100 33182 23214 33234
rect 23266 33182 23268 33234
rect 23100 33180 23268 33182
rect 22988 32562 23044 32574
rect 22988 32510 22990 32562
rect 23042 32510 23044 32562
rect 22876 31892 22932 31902
rect 22764 31890 22932 31892
rect 22764 31838 22878 31890
rect 22930 31838 22932 31890
rect 22764 31836 22932 31838
rect 22876 31826 22932 31836
rect 22988 31892 23044 32510
rect 22988 31826 23044 31836
rect 22652 31780 22708 31790
rect 22652 31686 22708 31724
rect 22428 31602 22484 31612
rect 22988 31554 23044 31566
rect 22988 31502 22990 31554
rect 23042 31502 23044 31554
rect 22988 31444 23044 31502
rect 22316 31388 23044 31444
rect 21756 31164 21924 31220
rect 21980 31332 22036 31342
rect 21756 30772 21812 31164
rect 21868 30996 21924 31006
rect 21980 30996 22036 31276
rect 21868 30994 22036 30996
rect 21868 30942 21870 30994
rect 21922 30942 22036 30994
rect 21868 30940 22036 30942
rect 21868 30930 21924 30940
rect 22092 30882 22148 30894
rect 22092 30830 22094 30882
rect 22146 30830 22148 30882
rect 21756 30716 21924 30772
rect 21644 30706 21700 30716
rect 21644 29988 21700 29998
rect 21644 29986 21812 29988
rect 21644 29934 21646 29986
rect 21698 29934 21812 29986
rect 21644 29932 21812 29934
rect 21644 29922 21700 29932
rect 21644 29316 21700 29326
rect 21644 29222 21700 29260
rect 21532 27794 21588 27804
rect 20412 27346 20468 27356
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 21756 24612 21812 29932
rect 21868 29652 21924 30716
rect 22092 30436 22148 30830
rect 22204 30436 22260 30446
rect 22092 30434 22260 30436
rect 22092 30382 22206 30434
rect 22258 30382 22260 30434
rect 22092 30380 22260 30382
rect 22204 30370 22260 30380
rect 21980 30098 22036 30110
rect 21980 30046 21982 30098
rect 22034 30046 22036 30098
rect 21980 29988 22036 30046
rect 22428 29988 22484 29998
rect 21980 29986 22484 29988
rect 21980 29934 22430 29986
rect 22482 29934 22484 29986
rect 21980 29932 22484 29934
rect 21980 29652 22036 29662
rect 21868 29650 22036 29652
rect 21868 29598 21982 29650
rect 22034 29598 22036 29650
rect 21868 29596 22036 29598
rect 21980 29202 22036 29596
rect 21980 29150 21982 29202
rect 22034 29150 22036 29202
rect 21980 29138 22036 29150
rect 21980 28756 22036 28766
rect 21980 28662 22036 28700
rect 21756 24546 21812 24556
rect 22428 24612 22484 29932
rect 22540 29650 22596 31388
rect 23100 31332 23156 33180
rect 23212 33170 23268 33180
rect 23324 33124 23380 33134
rect 23212 31668 23268 31678
rect 23212 31574 23268 31612
rect 23100 31266 23156 31276
rect 23212 31444 23268 31454
rect 22988 31108 23044 31118
rect 23212 31108 23268 31388
rect 23324 31218 23380 33068
rect 23436 33012 23492 33292
rect 23548 33346 23604 33358
rect 23548 33294 23550 33346
rect 23602 33294 23604 33346
rect 23548 33124 23604 33294
rect 23548 33058 23604 33068
rect 23436 32946 23492 32956
rect 23548 32788 23604 32798
rect 23324 31166 23326 31218
rect 23378 31166 23380 31218
rect 23324 31154 23380 31166
rect 23436 32676 23492 32686
rect 22988 31106 23268 31108
rect 22988 31054 22990 31106
rect 23042 31054 23268 31106
rect 22988 31052 23268 31054
rect 22988 31042 23044 31052
rect 22764 30996 22820 31006
rect 22764 30994 22932 30996
rect 22764 30942 22766 30994
rect 22818 30942 22932 30994
rect 22764 30940 22932 30942
rect 22764 30930 22820 30940
rect 22764 30434 22820 30446
rect 22764 30382 22766 30434
rect 22818 30382 22820 30434
rect 22540 29598 22542 29650
rect 22594 29598 22596 29650
rect 22540 29586 22596 29598
rect 22652 30212 22708 30222
rect 22540 29202 22596 29214
rect 22540 29150 22542 29202
rect 22594 29150 22596 29202
rect 22540 28754 22596 29150
rect 22540 28702 22542 28754
rect 22594 28702 22596 28754
rect 22540 28690 22596 28702
rect 22428 24546 22484 24556
rect 1820 10722 1876 10734
rect 1820 10670 1822 10722
rect 1874 10670 1876 10722
rect 1820 10164 1876 10670
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 1820 10098 1876 10108
rect 9100 9828 9156 9838
rect 9100 9714 9156 9772
rect 9100 9662 9102 9714
rect 9154 9662 9156 9714
rect 8764 9602 8820 9614
rect 8764 9550 8766 9602
rect 8818 9550 8820 9602
rect 1820 9154 1876 9166
rect 1820 9102 1822 9154
rect 1874 9102 1876 9154
rect 1820 8820 1876 9102
rect 1820 8754 1876 8764
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 1820 7586 1876 7598
rect 1820 7534 1822 7586
rect 1874 7534 1876 7586
rect 1820 6804 1876 7534
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 1820 6738 1876 6748
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 1820 4450 1876 4462
rect 1820 4398 1822 4450
rect 1874 4398 1876 4450
rect 1372 3556 1428 3566
rect 28 2324 84 2334
rect 28 800 84 2268
rect 1372 800 1428 3500
rect 1820 3444 1876 4398
rect 2492 4450 2548 4462
rect 2492 4398 2494 4450
rect 2546 4398 2548 4450
rect 2156 3556 2212 3566
rect 2156 3462 2212 3500
rect 1820 3378 1876 3388
rect 2492 2324 2548 4398
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 3052 3668 3108 3678
rect 3052 3554 3108 3612
rect 4284 3668 4340 3678
rect 4284 3574 4340 3612
rect 8764 3668 8820 9550
rect 9100 9604 9156 9662
rect 9100 9538 9156 9548
rect 9548 9604 9604 9614
rect 9548 9510 9604 9548
rect 12684 9604 12740 9614
rect 8764 3602 8820 3612
rect 3052 3502 3054 3554
rect 3106 3502 3108 3554
rect 3052 3490 3108 3502
rect 11900 3444 11956 3454
rect 12348 3444 12404 3454
rect 11900 3442 12404 3444
rect 11900 3390 11902 3442
rect 11954 3390 12350 3442
rect 12402 3390 12404 3442
rect 11900 3388 12404 3390
rect 11900 3378 11956 3388
rect 3612 3332 3668 3342
rect 2492 2258 2548 2268
rect 3388 3330 3668 3332
rect 3388 3278 3614 3330
rect 3666 3278 3668 3330
rect 3388 3276 3668 3278
rect 3388 800 3444 3276
rect 3612 3266 3668 3276
rect 4732 3332 4788 3342
rect 4732 800 4788 3276
rect 5740 3332 5796 3342
rect 5740 3238 5796 3276
rect 9660 3330 9716 3342
rect 9660 3278 9662 3330
rect 9714 3278 9716 3330
rect 8764 1762 8820 1774
rect 8764 1710 8766 1762
rect 8818 1710 8820 1762
rect 8764 800 8820 1710
rect 9660 1762 9716 3278
rect 9660 1710 9662 1762
rect 9714 1710 9716 1762
rect 9660 1698 9716 1710
rect 12124 800 12180 3388
rect 12348 3378 12404 3388
rect 12684 3330 12740 9548
rect 18620 3444 18676 3454
rect 19068 3444 19124 3454
rect 18620 3442 19124 3444
rect 18620 3390 18622 3442
rect 18674 3390 19070 3442
rect 19122 3390 19124 3442
rect 18620 3388 19124 3390
rect 18620 3378 18676 3388
rect 14364 3332 14420 3342
rect 15708 3332 15764 3342
rect 17724 3332 17780 3342
rect 12684 3278 12686 3330
rect 12738 3278 12740 3330
rect 12684 3266 12740 3278
rect 14140 3330 14420 3332
rect 14140 3278 14366 3330
rect 14418 3278 14420 3330
rect 14140 3276 14420 3278
rect 14140 800 14196 3276
rect 14364 3266 14420 3276
rect 15484 3330 15764 3332
rect 15484 3278 15710 3330
rect 15762 3278 15764 3330
rect 15484 3276 15764 3278
rect 15484 800 15540 3276
rect 15708 3266 15764 3276
rect 17500 3330 17780 3332
rect 17500 3278 17726 3330
rect 17778 3278 17780 3330
rect 17500 3276 17780 3278
rect 17500 800 17556 3276
rect 17724 3266 17780 3276
rect 18844 800 18900 3388
rect 19068 3378 19124 3388
rect 19404 3330 19460 11452
rect 19628 24500 19684 24510
rect 19628 11396 19684 24444
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 22652 18228 22708 30156
rect 22764 26180 22820 30382
rect 22876 29986 22932 30940
rect 22876 29934 22878 29986
rect 22930 29934 22932 29986
rect 22876 29204 22932 29934
rect 22988 30772 23044 30782
rect 22988 29650 23044 30716
rect 22988 29598 22990 29650
rect 23042 29598 23044 29650
rect 22988 29586 23044 29598
rect 23100 29652 23156 31052
rect 23436 30996 23492 32620
rect 23548 32674 23604 32732
rect 23548 32622 23550 32674
rect 23602 32622 23604 32674
rect 23548 32610 23604 32622
rect 23660 32450 23716 33404
rect 23996 33460 24052 35308
rect 23996 33394 24052 33404
rect 23884 33348 23940 33358
rect 23884 33254 23940 33292
rect 23660 32398 23662 32450
rect 23714 32398 23716 32450
rect 23660 32386 23716 32398
rect 23772 33124 23828 33134
rect 23772 32562 23828 33068
rect 24108 33124 24164 35980
rect 24220 35812 24276 35822
rect 24220 35028 24276 35756
rect 24220 34962 24276 34972
rect 24332 35588 24388 35598
rect 24220 34244 24276 34254
rect 24220 34130 24276 34188
rect 24220 34078 24222 34130
rect 24274 34078 24276 34130
rect 24220 34020 24276 34078
rect 24220 33954 24276 33964
rect 24108 33058 24164 33068
rect 24220 33796 24276 33806
rect 23772 32510 23774 32562
rect 23826 32510 23828 32562
rect 23772 32452 23828 32510
rect 23772 32386 23828 32396
rect 23884 32788 23940 32798
rect 23548 31668 23604 31678
rect 23548 31218 23604 31612
rect 23548 31166 23550 31218
rect 23602 31166 23604 31218
rect 23548 31154 23604 31166
rect 23772 31554 23828 31566
rect 23772 31502 23774 31554
rect 23826 31502 23828 31554
rect 23100 29586 23156 29596
rect 23212 30940 23492 30996
rect 22876 29138 22932 29148
rect 22988 28756 23044 28766
rect 22988 28662 23044 28700
rect 23212 28756 23268 30940
rect 23324 30770 23380 30782
rect 23324 30718 23326 30770
rect 23378 30718 23380 30770
rect 23324 29652 23380 30718
rect 23436 30434 23492 30446
rect 23436 30382 23438 30434
rect 23490 30382 23492 30434
rect 23436 30322 23492 30382
rect 23436 30270 23438 30322
rect 23490 30270 23492 30322
rect 23436 30258 23492 30270
rect 23436 29652 23492 29662
rect 23324 29650 23492 29652
rect 23324 29598 23438 29650
rect 23490 29598 23492 29650
rect 23324 29596 23492 29598
rect 23436 29586 23492 29596
rect 23212 28690 23268 28700
rect 22764 19908 22820 26124
rect 22764 19842 22820 19852
rect 22652 18162 22708 18172
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 23436 14868 23492 14878
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 23436 13188 23492 14812
rect 23436 13122 23492 13132
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 23772 11732 23828 31502
rect 23884 30660 23940 32732
rect 23996 32676 24052 32686
rect 23996 32582 24052 32620
rect 24220 32340 24276 33740
rect 24332 32900 24388 35532
rect 24444 34914 24500 36430
rect 24668 35588 24724 36988
rect 24780 35588 24836 35598
rect 24444 34862 24446 34914
rect 24498 34862 24500 34914
rect 24444 34850 24500 34862
rect 24556 35586 24836 35588
rect 24556 35534 24782 35586
rect 24834 35534 24836 35586
rect 24556 35532 24836 35534
rect 24444 34130 24500 34142
rect 24444 34078 24446 34130
rect 24498 34078 24500 34130
rect 24444 33124 24500 34078
rect 24556 33570 24612 35532
rect 24780 35522 24836 35532
rect 24892 35588 24948 35598
rect 24892 35494 24948 35532
rect 25116 34804 25172 37548
rect 25228 37156 25284 37996
rect 25228 37090 25284 37100
rect 25340 37604 25396 37614
rect 25340 37044 25396 37548
rect 25340 36978 25396 36988
rect 24668 34356 24724 34366
rect 24668 34262 24724 34300
rect 25004 34244 25060 34254
rect 24892 34130 24948 34142
rect 24892 34078 24894 34130
rect 24946 34078 24948 34130
rect 24780 34020 24836 34030
rect 24780 33926 24836 33964
rect 24556 33518 24558 33570
rect 24610 33518 24612 33570
rect 24556 33348 24612 33518
rect 24780 33684 24836 33694
rect 24780 33458 24836 33628
rect 24780 33406 24782 33458
rect 24834 33406 24836 33458
rect 24780 33394 24836 33406
rect 24892 33460 24948 34078
rect 25004 34020 25060 34188
rect 25004 33954 25060 33964
rect 24892 33394 24948 33404
rect 25004 33572 25060 33582
rect 24556 33282 24612 33292
rect 24780 33236 24836 33246
rect 24780 33142 24836 33180
rect 24444 33068 24724 33124
rect 24668 33012 24724 33068
rect 24668 32956 24836 33012
rect 24332 32844 24500 32900
rect 24444 32676 24500 32844
rect 24556 32676 24612 32686
rect 24444 32674 24612 32676
rect 24444 32622 24558 32674
rect 24610 32622 24612 32674
rect 24444 32620 24612 32622
rect 24556 32610 24612 32620
rect 24668 32676 24724 32686
rect 24220 32274 24276 32284
rect 24332 32452 24388 32462
rect 24108 31668 24164 31678
rect 23996 31666 24164 31668
rect 23996 31614 24110 31666
rect 24162 31614 24164 31666
rect 23996 31612 24164 31614
rect 23996 31108 24052 31612
rect 24108 31602 24164 31612
rect 23996 31014 24052 31052
rect 23884 30594 23940 30604
rect 23996 30324 24052 30334
rect 23884 30212 23940 30222
rect 23884 30118 23940 30156
rect 23884 29652 23940 29662
rect 23996 29652 24052 30268
rect 24332 30322 24388 32396
rect 24668 31890 24724 32620
rect 24668 31838 24670 31890
rect 24722 31838 24724 31890
rect 24668 31826 24724 31838
rect 24444 30884 24500 30894
rect 24444 30436 24500 30828
rect 24444 30370 24500 30380
rect 24332 30270 24334 30322
rect 24386 30270 24388 30322
rect 24332 30258 24388 30270
rect 24780 29988 24836 32956
rect 24892 32788 24948 32798
rect 24892 32674 24948 32732
rect 24892 32622 24894 32674
rect 24946 32622 24948 32674
rect 24892 32610 24948 32622
rect 25004 32564 25060 33516
rect 24892 31220 24948 31230
rect 25004 31220 25060 32508
rect 24892 31218 25060 31220
rect 24892 31166 24894 31218
rect 24946 31166 25060 31218
rect 24892 31164 25060 31166
rect 24892 31154 24948 31164
rect 25116 30324 25172 34748
rect 25228 36708 25284 36718
rect 25228 35700 25284 36652
rect 25340 36484 25396 36494
rect 25340 36390 25396 36428
rect 25228 34914 25284 35644
rect 25228 34862 25230 34914
rect 25282 34862 25284 34914
rect 25228 34692 25284 34862
rect 25452 35252 25508 41244
rect 25788 40402 25844 40414
rect 25788 40350 25790 40402
rect 25842 40350 25844 40402
rect 25788 40180 25844 40350
rect 25788 40114 25844 40124
rect 25788 38948 25844 38958
rect 25676 38836 25732 38846
rect 25676 38722 25732 38780
rect 25676 38670 25678 38722
rect 25730 38670 25732 38722
rect 25676 38658 25732 38670
rect 25676 37156 25732 37166
rect 25452 35138 25508 35196
rect 25452 35086 25454 35138
rect 25506 35086 25508 35138
rect 25228 34626 25284 34636
rect 25340 34690 25396 34702
rect 25340 34638 25342 34690
rect 25394 34638 25396 34690
rect 25228 32900 25284 32910
rect 25228 31890 25284 32844
rect 25228 31838 25230 31890
rect 25282 31838 25284 31890
rect 25228 31826 25284 31838
rect 25340 31780 25396 34638
rect 25452 34132 25508 35086
rect 25452 34066 25508 34076
rect 25564 37154 25732 37156
rect 25564 37102 25678 37154
rect 25730 37102 25732 37154
rect 25564 37100 25732 37102
rect 25564 33348 25620 37100
rect 25676 37090 25732 37100
rect 25676 35700 25732 35710
rect 25676 35606 25732 35644
rect 25676 35140 25732 35150
rect 25788 35140 25844 38892
rect 25900 38500 25956 38510
rect 25900 37938 25956 38444
rect 25900 37886 25902 37938
rect 25954 37886 25956 37938
rect 25900 37828 25956 37886
rect 25900 37762 25956 37772
rect 25900 37380 25956 37390
rect 25900 37286 25956 37324
rect 26012 37156 26068 45166
rect 26124 42308 26180 45836
rect 26124 42242 26180 42252
rect 26348 38724 26404 45950
rect 26572 45106 26628 47964
rect 26908 45780 26964 49200
rect 27020 48802 27076 48814
rect 27020 48750 27022 48802
rect 27074 48750 27076 48802
rect 27020 48692 27076 48750
rect 27020 48626 27076 48636
rect 30156 48580 30212 48590
rect 28812 48356 28868 48366
rect 27020 48020 27076 48030
rect 27020 47794 27076 47964
rect 27020 47742 27022 47794
rect 27074 47742 27076 47794
rect 27020 47730 27076 47742
rect 27804 47684 27860 47694
rect 27244 47572 27300 47582
rect 26908 45714 26964 45724
rect 27020 46900 27076 46910
rect 26572 45054 26574 45106
rect 26626 45054 26628 45106
rect 26572 45042 26628 45054
rect 27020 45332 27076 46844
rect 26908 44882 26964 44894
rect 26908 44830 26910 44882
rect 26962 44830 26964 44882
rect 26684 44772 26740 44782
rect 26460 41860 26516 41870
rect 26460 41858 26628 41860
rect 26460 41806 26462 41858
rect 26514 41806 26628 41858
rect 26460 41804 26628 41806
rect 26460 41794 26516 41804
rect 26460 41188 26516 41198
rect 26460 40852 26516 41132
rect 26460 40514 26516 40796
rect 26460 40462 26462 40514
rect 26514 40462 26516 40514
rect 26460 40450 26516 40462
rect 26348 38658 26404 38668
rect 26460 40292 26516 40302
rect 26012 37090 26068 37100
rect 26236 38164 26292 38174
rect 26124 37044 26180 37054
rect 26012 36708 26068 36718
rect 26012 36594 26068 36652
rect 26124 36706 26180 36988
rect 26124 36654 26126 36706
rect 26178 36654 26180 36706
rect 26124 36642 26180 36654
rect 26012 36542 26014 36594
rect 26066 36542 26068 36594
rect 26012 36530 26068 36542
rect 26012 36372 26068 36382
rect 25900 36148 25956 36158
rect 25900 35810 25956 36092
rect 25900 35758 25902 35810
rect 25954 35758 25956 35810
rect 25900 35746 25956 35758
rect 25676 35138 25956 35140
rect 25676 35086 25678 35138
rect 25730 35086 25956 35138
rect 25676 35084 25956 35086
rect 25676 35074 25732 35084
rect 25788 34914 25844 34926
rect 25788 34862 25790 34914
rect 25842 34862 25844 34914
rect 25788 34804 25844 34862
rect 25788 34738 25844 34748
rect 25676 34244 25732 34254
rect 25676 34150 25732 34188
rect 25676 33348 25732 33358
rect 25564 33346 25732 33348
rect 25564 33294 25678 33346
rect 25730 33294 25732 33346
rect 25564 33292 25732 33294
rect 25676 33282 25732 33292
rect 25452 33236 25508 33246
rect 25452 33142 25508 33180
rect 25340 31714 25396 31724
rect 25564 33012 25620 33022
rect 25564 31220 25620 32956
rect 25676 32788 25732 32798
rect 25676 32694 25732 32732
rect 25676 31892 25732 31902
rect 25676 31798 25732 31836
rect 25900 31780 25956 35084
rect 26012 34468 26068 36316
rect 26124 35476 26180 35486
rect 26124 35382 26180 35420
rect 26012 34402 26068 34412
rect 26012 34244 26068 34254
rect 26012 34242 26180 34244
rect 26012 34190 26014 34242
rect 26066 34190 26180 34242
rect 26012 34188 26180 34190
rect 26012 34178 26068 34188
rect 26012 33124 26068 33134
rect 26012 32786 26068 33068
rect 26012 32734 26014 32786
rect 26066 32734 26068 32786
rect 26012 32676 26068 32734
rect 26012 32610 26068 32620
rect 26124 31780 26180 34188
rect 26236 33460 26292 38108
rect 26348 36596 26404 36606
rect 26348 35698 26404 36540
rect 26460 35922 26516 40236
rect 26572 38668 26628 41804
rect 26684 41186 26740 44716
rect 26908 41972 26964 44830
rect 26908 41906 26964 41916
rect 26908 41300 26964 41310
rect 26908 41206 26964 41244
rect 26684 41134 26686 41186
rect 26738 41134 26740 41186
rect 26684 39620 26740 41134
rect 27020 41074 27076 45276
rect 27020 41022 27022 41074
rect 27074 41022 27076 41074
rect 27020 41010 27076 41022
rect 27132 45444 27188 45454
rect 26684 39554 26740 39564
rect 27132 39732 27188 45388
rect 27244 42866 27300 47516
rect 27804 47124 27860 47628
rect 27580 46564 27636 46574
rect 27356 45892 27412 45902
rect 27356 45778 27412 45836
rect 27356 45726 27358 45778
rect 27410 45726 27412 45778
rect 27356 45714 27412 45726
rect 27468 45778 27524 45790
rect 27468 45726 27470 45778
rect 27522 45726 27524 45778
rect 27468 45444 27524 45726
rect 27580 45778 27636 46508
rect 27692 46562 27748 46574
rect 27692 46510 27694 46562
rect 27746 46510 27748 46562
rect 27692 46116 27748 46510
rect 27692 46050 27748 46060
rect 27804 45890 27860 47068
rect 28364 46228 28420 46238
rect 28028 46116 28084 46126
rect 27804 45838 27806 45890
rect 27858 45838 27860 45890
rect 27804 45826 27860 45838
rect 27916 46004 27972 46014
rect 27580 45726 27582 45778
rect 27634 45726 27636 45778
rect 27580 45714 27636 45726
rect 27692 45668 27748 45678
rect 27692 45574 27748 45612
rect 27468 45378 27524 45388
rect 27804 45556 27860 45566
rect 27580 44996 27636 45006
rect 27580 44902 27636 44940
rect 27244 42814 27246 42866
rect 27298 42814 27300 42866
rect 27244 39956 27300 42814
rect 27692 43764 27748 43774
rect 27244 39890 27300 39900
rect 27356 41636 27412 41646
rect 26908 38724 26964 38734
rect 26572 38612 26740 38668
rect 26460 35870 26462 35922
rect 26514 35870 26516 35922
rect 26460 35858 26516 35870
rect 26348 35646 26350 35698
rect 26402 35646 26404 35698
rect 26348 35634 26404 35646
rect 26572 35698 26628 35710
rect 26572 35646 26574 35698
rect 26626 35646 26628 35698
rect 26572 35364 26628 35646
rect 26572 35298 26628 35308
rect 26460 34690 26516 34702
rect 26460 34638 26462 34690
rect 26514 34638 26516 34690
rect 26348 33460 26404 33470
rect 26236 33458 26404 33460
rect 26236 33406 26350 33458
rect 26402 33406 26404 33458
rect 26236 33404 26404 33406
rect 26348 33394 26404 33404
rect 26460 33348 26516 34638
rect 26572 34356 26628 34366
rect 26684 34356 26740 38612
rect 26796 36372 26852 36382
rect 26796 36278 26852 36316
rect 26572 34354 26740 34356
rect 26572 34302 26574 34354
rect 26626 34302 26740 34354
rect 26572 34300 26740 34302
rect 26796 34914 26852 34926
rect 26796 34862 26798 34914
rect 26850 34862 26852 34914
rect 26572 34290 26628 34300
rect 26796 34020 26852 34862
rect 26908 34356 26964 38668
rect 27132 38164 27188 39676
rect 27244 39508 27300 39518
rect 27244 39060 27300 39452
rect 27244 38994 27300 39004
rect 27132 38108 27300 38164
rect 27132 37828 27188 37838
rect 27020 37268 27076 37278
rect 27020 37174 27076 37212
rect 27132 37156 27188 37772
rect 27244 37378 27300 38108
rect 27244 37326 27246 37378
rect 27298 37326 27300 37378
rect 27244 37314 27300 37326
rect 27132 37100 27300 37156
rect 27132 36484 27188 36494
rect 27020 36428 27132 36484
rect 27020 35924 27076 36428
rect 27132 36390 27188 36428
rect 27244 36482 27300 37100
rect 27244 36430 27246 36482
rect 27298 36430 27300 36482
rect 27244 36372 27300 36430
rect 27244 36306 27300 36316
rect 27020 35858 27076 35868
rect 27132 35924 27188 35934
rect 27356 35924 27412 41580
rect 27692 41186 27748 43708
rect 27804 43650 27860 45500
rect 27916 44436 27972 45948
rect 28028 45556 28084 46060
rect 28364 46114 28420 46172
rect 28364 46062 28366 46114
rect 28418 46062 28420 46114
rect 28364 46050 28420 46062
rect 28476 45780 28532 45790
rect 28028 45490 28084 45500
rect 28252 45778 28532 45780
rect 28252 45726 28478 45778
rect 28530 45726 28532 45778
rect 28252 45724 28532 45726
rect 28028 45220 28084 45230
rect 28028 44660 28084 45164
rect 28140 45108 28196 45118
rect 28140 45014 28196 45052
rect 28028 44594 28084 44604
rect 28028 44436 28084 44446
rect 27916 44434 28084 44436
rect 27916 44382 28030 44434
rect 28082 44382 28084 44434
rect 27916 44380 28084 44382
rect 27804 43598 27806 43650
rect 27858 43598 27860 43650
rect 27804 43316 27860 43598
rect 27804 43250 27860 43260
rect 27692 41134 27694 41186
rect 27746 41134 27748 41186
rect 27692 41122 27748 41134
rect 27916 42756 27972 42766
rect 27916 41188 27972 42700
rect 27916 40180 27972 41132
rect 28028 40516 28084 44380
rect 28252 41636 28308 45724
rect 28476 45714 28532 45724
rect 28700 45444 28756 45454
rect 28364 45106 28420 45118
rect 28364 45054 28366 45106
rect 28418 45054 28420 45106
rect 28364 44996 28420 45054
rect 28364 44212 28420 44940
rect 28700 44546 28756 45388
rect 28700 44494 28702 44546
rect 28754 44494 28756 44546
rect 28700 44482 28756 44494
rect 28812 44436 28868 48300
rect 29372 48356 29428 48366
rect 28924 47796 28980 47806
rect 28924 45218 28980 47740
rect 29260 45666 29316 45678
rect 29260 45614 29262 45666
rect 29314 45614 29316 45666
rect 29260 45556 29316 45614
rect 29260 45490 29316 45500
rect 29372 45332 29428 48300
rect 29820 47908 29876 47918
rect 29708 47852 29820 47908
rect 28924 45166 28926 45218
rect 28978 45166 28980 45218
rect 28924 45154 28980 45166
rect 29260 45276 29428 45332
rect 29484 47684 29540 47694
rect 29260 45218 29316 45276
rect 29260 45166 29262 45218
rect 29314 45166 29316 45218
rect 29260 45154 29316 45166
rect 29372 45106 29428 45118
rect 29372 45054 29374 45106
rect 29426 45054 29428 45106
rect 29036 44994 29092 45006
rect 29036 44942 29038 44994
rect 29090 44942 29092 44994
rect 28812 44380 28980 44436
rect 28364 43708 28420 44156
rect 28700 44324 28756 44334
rect 28700 44210 28756 44268
rect 28700 44158 28702 44210
rect 28754 44158 28756 44210
rect 28700 44146 28756 44158
rect 28812 44212 28868 44222
rect 28364 43652 28756 43708
rect 28476 43538 28532 43550
rect 28476 43486 28478 43538
rect 28530 43486 28532 43538
rect 28476 42756 28532 43486
rect 28700 42978 28756 43652
rect 28700 42926 28702 42978
rect 28754 42926 28756 42978
rect 28700 42914 28756 42926
rect 28476 42690 28532 42700
rect 28588 42756 28644 42766
rect 28812 42756 28868 44156
rect 28924 43316 28980 44380
rect 29036 43764 29092 44942
rect 29372 44884 29428 45054
rect 29372 44818 29428 44828
rect 29484 44324 29540 47628
rect 29596 45668 29652 45678
rect 29596 45574 29652 45612
rect 29708 44996 29764 47852
rect 29820 47842 29876 47852
rect 30156 47796 30212 48524
rect 30156 47730 30212 47740
rect 30604 48468 30660 48478
rect 30604 47796 30660 48412
rect 30380 47236 30436 47246
rect 29820 46562 29876 46574
rect 29820 46510 29822 46562
rect 29874 46510 29876 46562
rect 29820 45556 29876 46510
rect 30156 45780 30212 45790
rect 30156 45686 30212 45724
rect 29820 45490 29876 45500
rect 30380 45220 30436 47180
rect 30604 46340 30660 47740
rect 30828 48468 30884 48478
rect 30604 46274 30660 46284
rect 30716 47460 30772 47470
rect 30268 45218 30436 45220
rect 30268 45166 30382 45218
rect 30434 45166 30436 45218
rect 30268 45164 30436 45166
rect 30044 45108 30100 45146
rect 30044 45042 30100 45052
rect 29708 44930 29764 44940
rect 30156 44996 30212 45006
rect 30044 44884 30100 44894
rect 29932 44882 30100 44884
rect 29932 44830 30046 44882
rect 30098 44830 30100 44882
rect 29932 44828 30100 44830
rect 29708 44324 29764 44334
rect 29484 44258 29540 44268
rect 29596 44268 29708 44324
rect 29596 44100 29652 44268
rect 29708 44258 29764 44268
rect 29820 44324 29876 44334
rect 29932 44324 29988 44828
rect 30044 44818 30100 44828
rect 29820 44322 29988 44324
rect 29820 44270 29822 44322
rect 29874 44270 29988 44322
rect 29820 44268 29988 44270
rect 29820 44258 29876 44268
rect 29036 43698 29092 43708
rect 29372 44098 29652 44100
rect 29372 44046 29598 44098
rect 29650 44046 29652 44098
rect 29372 44044 29652 44046
rect 29036 43428 29092 43438
rect 29036 43334 29092 43372
rect 28924 43250 28980 43260
rect 29372 42868 29428 44044
rect 29596 44034 29652 44044
rect 29708 44098 29764 44110
rect 29708 44046 29710 44098
rect 29762 44046 29764 44098
rect 29484 43876 29540 43886
rect 29484 43538 29540 43820
rect 29708 43708 29764 44046
rect 30044 44100 30100 44110
rect 30044 44006 30100 44044
rect 29484 43486 29486 43538
rect 29538 43486 29540 43538
rect 29484 43474 29540 43486
rect 29596 43652 29764 43708
rect 30044 43652 30100 43662
rect 29372 42802 29428 42812
rect 28588 42754 28868 42756
rect 28588 42702 28590 42754
rect 28642 42702 28868 42754
rect 28588 42700 28868 42702
rect 28588 42690 28644 42700
rect 28700 42530 28756 42542
rect 28700 42478 28702 42530
rect 28754 42478 28756 42530
rect 28588 42308 28644 42318
rect 28588 41858 28644 42252
rect 28700 42084 28756 42478
rect 28700 42018 28756 42028
rect 28588 41806 28590 41858
rect 28642 41806 28644 41858
rect 28588 41794 28644 41806
rect 28588 41636 28644 41646
rect 28252 41580 28532 41636
rect 28028 40450 28084 40460
rect 28252 41412 28308 41422
rect 28252 41186 28308 41356
rect 28252 41134 28254 41186
rect 28306 41134 28308 41186
rect 27916 39618 27972 40124
rect 27916 39566 27918 39618
rect 27970 39566 27972 39618
rect 27468 39396 27524 39406
rect 27468 37828 27524 39340
rect 27804 38948 27860 38958
rect 27804 38854 27860 38892
rect 27916 38836 27972 39566
rect 27916 38770 27972 38780
rect 28028 39956 28084 39966
rect 27468 37762 27524 37772
rect 28028 38162 28084 39900
rect 28028 38110 28030 38162
rect 28082 38110 28084 38162
rect 27804 37380 27860 37390
rect 27692 36820 27748 36830
rect 27580 36764 27692 36820
rect 27468 36596 27524 36606
rect 27580 36596 27636 36764
rect 27692 36754 27748 36764
rect 27468 36594 27636 36596
rect 27468 36542 27470 36594
rect 27522 36542 27636 36594
rect 27468 36540 27636 36542
rect 27468 36530 27524 36540
rect 27692 36370 27748 36382
rect 27692 36318 27694 36370
rect 27746 36318 27748 36370
rect 27132 35922 27412 35924
rect 27132 35870 27134 35922
rect 27186 35870 27412 35922
rect 27132 35868 27412 35870
rect 27468 36036 27524 36046
rect 27132 35858 27188 35868
rect 27468 35812 27524 35980
rect 27692 35924 27748 36318
rect 27804 36258 27860 37324
rect 27804 36206 27806 36258
rect 27858 36206 27860 36258
rect 27804 36194 27860 36206
rect 28028 36036 28084 38110
rect 28028 35970 28084 35980
rect 28140 39620 28196 39630
rect 27692 35858 27748 35868
rect 27244 35756 27524 35812
rect 28140 35812 28196 39564
rect 28252 39284 28308 41134
rect 28476 39620 28532 41580
rect 28588 40290 28644 41580
rect 28812 41524 28868 42700
rect 28812 41458 28868 41468
rect 28924 42756 28980 42766
rect 28700 40964 28756 40974
rect 28700 40962 28868 40964
rect 28700 40910 28702 40962
rect 28754 40910 28868 40962
rect 28700 40908 28868 40910
rect 28700 40898 28756 40908
rect 28588 40238 28590 40290
rect 28642 40238 28644 40290
rect 28588 40226 28644 40238
rect 28700 40068 28756 40078
rect 28700 39842 28756 40012
rect 28700 39790 28702 39842
rect 28754 39790 28756 39842
rect 28700 39778 28756 39790
rect 28588 39620 28644 39630
rect 28532 39618 28644 39620
rect 28532 39566 28590 39618
rect 28642 39566 28644 39618
rect 28532 39564 28644 39566
rect 28476 39488 28532 39564
rect 28588 39554 28644 39564
rect 28700 39396 28756 39406
rect 28700 39302 28756 39340
rect 28252 39228 28420 39284
rect 28364 36932 28420 39228
rect 28812 39172 28868 40908
rect 28924 39508 28980 42700
rect 29484 42532 29540 42542
rect 29372 42530 29540 42532
rect 29372 42478 29486 42530
rect 29538 42478 29540 42530
rect 29372 42476 29540 42478
rect 29148 41524 29204 41534
rect 29372 41524 29428 42476
rect 29484 42466 29540 42476
rect 29148 40516 29204 41468
rect 29260 41468 29428 41524
rect 29484 41972 29540 41982
rect 29260 40740 29316 41468
rect 29260 40674 29316 40684
rect 29372 41300 29428 41310
rect 29372 40628 29428 41244
rect 29260 40516 29316 40526
rect 29148 40514 29316 40516
rect 29148 40462 29262 40514
rect 29314 40462 29316 40514
rect 29148 40460 29316 40462
rect 29260 40450 29316 40460
rect 29372 40402 29428 40572
rect 29372 40350 29374 40402
rect 29426 40350 29428 40402
rect 29372 40338 29428 40350
rect 29484 40740 29540 41916
rect 29596 41524 29652 43652
rect 29708 43538 29764 43550
rect 29708 43486 29710 43538
rect 29762 43486 29764 43538
rect 29708 42756 29764 43486
rect 29820 43538 29876 43550
rect 29820 43486 29822 43538
rect 29874 43486 29876 43538
rect 29820 43428 29876 43486
rect 30044 43538 30100 43596
rect 30044 43486 30046 43538
rect 30098 43486 30100 43538
rect 30044 43474 30100 43486
rect 29820 43362 29876 43372
rect 29932 43316 29988 43326
rect 29932 42978 29988 43260
rect 30156 43204 30212 44940
rect 29932 42926 29934 42978
rect 29986 42926 29988 42978
rect 29932 42914 29988 42926
rect 30044 43148 30212 43204
rect 29708 42690 29764 42700
rect 29820 42868 29876 42878
rect 29820 42532 29876 42812
rect 30044 42532 30100 43148
rect 30156 42868 30212 42878
rect 30156 42774 30212 42812
rect 30044 42476 30212 42532
rect 29820 42466 29876 42476
rect 29932 42084 29988 42094
rect 29820 41972 29876 41982
rect 29596 41468 29764 41524
rect 29596 41300 29652 41310
rect 29596 41206 29652 41244
rect 29484 39844 29540 40684
rect 29708 40292 29764 41468
rect 29708 40226 29764 40236
rect 29820 40180 29876 41916
rect 29932 41746 29988 42028
rect 29932 41694 29934 41746
rect 29986 41694 29988 41746
rect 29932 41682 29988 41694
rect 30044 41970 30100 41982
rect 30044 41918 30046 41970
rect 30098 41918 30100 41970
rect 30044 41524 30100 41918
rect 30044 41458 30100 41468
rect 29820 40114 29876 40124
rect 29932 41076 29988 41086
rect 29820 39956 29876 39966
rect 29596 39844 29652 39854
rect 29484 39842 29652 39844
rect 29484 39790 29598 39842
rect 29650 39790 29652 39842
rect 29484 39788 29652 39790
rect 29596 39778 29652 39788
rect 29820 39842 29876 39900
rect 29820 39790 29822 39842
rect 29874 39790 29876 39842
rect 29820 39778 29876 39790
rect 28924 39452 29092 39508
rect 28700 39116 28868 39172
rect 28476 38836 28532 38846
rect 28476 38742 28532 38780
rect 28700 38500 28756 39116
rect 28700 38434 28756 38444
rect 28812 38948 28868 38958
rect 28812 38164 28868 38892
rect 28476 38108 28868 38164
rect 28476 37044 28532 38108
rect 28924 38052 28980 38062
rect 28812 37996 28924 38052
rect 28588 37938 28644 37950
rect 28588 37886 28590 37938
rect 28642 37886 28644 37938
rect 28588 37604 28644 37886
rect 28700 37828 28756 37838
rect 28700 37734 28756 37772
rect 28812 37604 28868 37996
rect 28924 37986 28980 37996
rect 29036 37940 29092 39452
rect 29372 39396 29428 39406
rect 29260 38948 29316 38958
rect 29372 38948 29428 39340
rect 29820 39284 29876 39294
rect 29484 38948 29540 38958
rect 29372 38946 29540 38948
rect 29372 38894 29486 38946
rect 29538 38894 29540 38946
rect 29372 38892 29540 38894
rect 29260 38854 29316 38892
rect 29484 38882 29540 38892
rect 29708 38948 29764 38958
rect 29820 38948 29876 39228
rect 29708 38946 29876 38948
rect 29708 38894 29710 38946
rect 29762 38894 29876 38946
rect 29708 38892 29876 38894
rect 29148 38722 29204 38734
rect 29148 38670 29150 38722
rect 29202 38670 29204 38722
rect 29148 38164 29204 38670
rect 29708 38276 29764 38892
rect 29932 38388 29988 41020
rect 30044 40516 30100 40526
rect 30044 40402 30100 40460
rect 30044 40350 30046 40402
rect 30098 40350 30100 40402
rect 30044 40338 30100 40350
rect 30156 39618 30212 42476
rect 30268 40964 30324 45164
rect 30380 45154 30436 45164
rect 30716 44322 30772 47404
rect 30828 47236 30884 48412
rect 30828 47170 30884 47180
rect 30940 45780 30996 49200
rect 30940 45714 30996 45724
rect 31276 48692 31332 48702
rect 31164 45668 31220 45678
rect 31052 45666 31220 45668
rect 31052 45614 31166 45666
rect 31218 45614 31220 45666
rect 31052 45612 31220 45614
rect 30716 44270 30718 44322
rect 30770 44270 30772 44322
rect 30716 44258 30772 44270
rect 30828 45108 30884 45118
rect 30828 44100 30884 45052
rect 31052 44996 31108 45612
rect 31164 45602 31220 45612
rect 31052 44902 31108 44940
rect 30940 44882 30996 44894
rect 30940 44830 30942 44882
rect 30994 44830 30996 44882
rect 30940 44660 30996 44830
rect 30940 44594 30996 44604
rect 31052 44772 31108 44782
rect 31052 44322 31108 44716
rect 31164 44548 31220 44558
rect 31276 44548 31332 48636
rect 31836 48244 31892 48254
rect 31836 47460 31892 48188
rect 31836 47394 31892 47404
rect 31948 47236 32004 49196
rect 31948 47170 32004 47180
rect 31948 46562 32004 46574
rect 31948 46510 31950 46562
rect 32002 46510 32004 46562
rect 31500 45780 31556 45790
rect 31500 45686 31556 45724
rect 31500 45332 31556 45342
rect 31948 45332 32004 46510
rect 32060 45778 32116 49868
rect 32508 49812 32564 49822
rect 32256 49200 32368 49800
rect 32284 46786 32340 49200
rect 32284 46734 32286 46786
rect 32338 46734 32340 46786
rect 32284 46722 32340 46734
rect 32396 48132 32452 48142
rect 32284 46564 32340 46574
rect 32060 45726 32062 45778
rect 32114 45726 32116 45778
rect 32060 45714 32116 45726
rect 32172 45892 32228 45902
rect 32172 45668 32228 45836
rect 32060 45332 32116 45342
rect 31948 45330 32116 45332
rect 31948 45278 32062 45330
rect 32114 45278 32116 45330
rect 31948 45276 32116 45278
rect 31500 45238 31556 45276
rect 32060 45266 32116 45276
rect 31948 44882 32004 44894
rect 31948 44830 31950 44882
rect 32002 44830 32004 44882
rect 31220 44492 31332 44548
rect 31836 44548 31892 44558
rect 31164 44434 31220 44492
rect 31164 44382 31166 44434
rect 31218 44382 31220 44434
rect 31164 44370 31220 44382
rect 31052 44270 31054 44322
rect 31106 44270 31108 44322
rect 31052 44258 31108 44270
rect 31836 44322 31892 44492
rect 31836 44270 31838 44322
rect 31890 44270 31892 44322
rect 31836 44258 31892 44270
rect 30828 44044 31108 44100
rect 30380 43988 30436 43998
rect 30380 42978 30436 43932
rect 30380 42926 30382 42978
rect 30434 42926 30436 42978
rect 30380 42914 30436 42926
rect 30492 43764 30548 43774
rect 30380 42756 30436 42766
rect 30380 42532 30436 42700
rect 30380 42466 30436 42476
rect 30380 41970 30436 41982
rect 30380 41918 30382 41970
rect 30434 41918 30436 41970
rect 30380 41748 30436 41918
rect 30492 41858 30548 43708
rect 31052 43762 31108 44044
rect 31052 43710 31054 43762
rect 31106 43710 31108 43762
rect 31052 43698 31108 43710
rect 31276 44098 31332 44110
rect 31276 44046 31278 44098
rect 31330 44046 31332 44098
rect 31276 43708 31332 44046
rect 31724 44100 31780 44110
rect 31724 43762 31780 44044
rect 31724 43710 31726 43762
rect 31778 43710 31780 43762
rect 30604 43652 30660 43662
rect 31276 43652 31668 43708
rect 31724 43698 31780 43710
rect 30604 42866 30660 43596
rect 30604 42814 30606 42866
rect 30658 42814 30660 42866
rect 30604 42802 30660 42814
rect 30716 43538 30772 43550
rect 30716 43486 30718 43538
rect 30770 43486 30772 43538
rect 30716 42196 30772 43486
rect 30492 41806 30494 41858
rect 30546 41806 30548 41858
rect 30492 41794 30548 41806
rect 30604 42140 30772 42196
rect 30828 43538 30884 43550
rect 30828 43486 30830 43538
rect 30882 43486 30884 43538
rect 30380 41682 30436 41692
rect 30268 40898 30324 40908
rect 30380 41076 30436 41086
rect 30268 40514 30324 40526
rect 30268 40462 30270 40514
rect 30322 40462 30324 40514
rect 30268 39844 30324 40462
rect 30268 39778 30324 39788
rect 30156 39566 30158 39618
rect 30210 39566 30212 39618
rect 30156 39554 30212 39566
rect 30268 39620 30324 39630
rect 30380 39620 30436 41020
rect 30604 39732 30660 42140
rect 30716 41972 30772 41982
rect 30716 41878 30772 41916
rect 30604 39666 30660 39676
rect 30828 41300 30884 43486
rect 30940 43540 30996 43578
rect 30940 43474 30996 43484
rect 31276 43540 31332 43550
rect 31276 43446 31332 43484
rect 31500 43540 31556 43550
rect 31500 43316 31556 43484
rect 31276 43260 31556 43316
rect 31276 42756 31332 43260
rect 31612 42868 31668 43652
rect 31836 43650 31892 43662
rect 31836 43598 31838 43650
rect 31890 43598 31892 43650
rect 31836 43540 31892 43598
rect 31612 42812 31780 42868
rect 31276 42690 31332 42700
rect 31500 42756 31556 42766
rect 31388 42644 31444 42654
rect 31164 42530 31220 42542
rect 31164 42478 31166 42530
rect 31218 42478 31220 42530
rect 31164 41860 31220 42478
rect 31164 41794 31220 41804
rect 31276 42530 31332 42542
rect 31276 42478 31278 42530
rect 31330 42478 31332 42530
rect 30268 39618 30436 39620
rect 30268 39566 30270 39618
rect 30322 39566 30436 39618
rect 30268 39564 30436 39566
rect 30268 39554 30324 39564
rect 30380 39394 30436 39406
rect 30380 39342 30382 39394
rect 30434 39342 30436 39394
rect 30380 39172 30436 39342
rect 30492 39396 30548 39406
rect 30492 39302 30548 39340
rect 30828 39172 30884 41244
rect 30940 40404 30996 40414
rect 30940 40310 30996 40348
rect 31164 39732 31220 39742
rect 31164 39638 31220 39676
rect 31276 39396 31332 42478
rect 31388 41748 31444 42588
rect 31500 42642 31556 42700
rect 31500 42590 31502 42642
rect 31554 42590 31556 42642
rect 31500 42578 31556 42590
rect 31612 42644 31668 42654
rect 31612 42550 31668 42588
rect 31724 42420 31780 42812
rect 31836 42644 31892 43484
rect 31836 42578 31892 42588
rect 31388 41682 31444 41692
rect 31500 42364 31780 42420
rect 31500 41412 31556 42364
rect 31948 42308 32004 44830
rect 32172 44772 32228 45612
rect 32060 44716 32228 44772
rect 32060 43650 32116 44716
rect 32172 44212 32228 44222
rect 32284 44212 32340 46508
rect 32172 44210 32340 44212
rect 32172 44158 32174 44210
rect 32226 44158 32340 44210
rect 32172 44156 32340 44158
rect 32396 45330 32452 48076
rect 32396 45278 32398 45330
rect 32450 45278 32452 45330
rect 32172 44146 32228 44156
rect 32396 43764 32452 45278
rect 32396 43698 32452 43708
rect 32060 43598 32062 43650
rect 32114 43598 32116 43650
rect 32060 43586 32116 43598
rect 32396 43540 32452 43550
rect 32508 43540 32564 49756
rect 34272 49200 34384 49800
rect 34972 49588 35028 49598
rect 35028 49532 35140 49588
rect 34972 49522 35028 49532
rect 34300 47348 34356 47358
rect 33068 47236 33124 47246
rect 32844 44994 32900 45006
rect 32844 44942 32846 44994
rect 32898 44942 32900 44994
rect 32844 44882 32900 44942
rect 32844 44830 32846 44882
rect 32898 44830 32900 44882
rect 32844 44818 32900 44830
rect 33068 44434 33124 47180
rect 33404 46786 33460 46798
rect 33404 46734 33406 46786
rect 33458 46734 33460 46786
rect 33404 46002 33460 46734
rect 33404 45950 33406 46002
rect 33458 45950 33460 46002
rect 33404 45938 33460 45950
rect 33628 46116 33684 46126
rect 33068 44382 33070 44434
rect 33122 44382 33124 44434
rect 33068 44370 33124 44382
rect 33628 45108 33684 46060
rect 32732 44100 32788 44110
rect 32732 44006 32788 44044
rect 33516 44098 33572 44110
rect 33516 44046 33518 44098
rect 33570 44046 33572 44098
rect 33516 43988 33572 44046
rect 32396 43538 32508 43540
rect 32396 43486 32398 43538
rect 32450 43486 32508 43538
rect 32396 43484 32508 43486
rect 32396 43474 32452 43484
rect 32508 43408 32564 43484
rect 33068 43932 33572 43988
rect 32732 43426 32788 43438
rect 32732 43374 32734 43426
rect 32786 43374 32788 43426
rect 31948 42242 32004 42252
rect 32396 43204 32452 43214
rect 31948 42084 32004 42094
rect 31948 41990 32004 42028
rect 32172 42084 32228 42094
rect 31836 41972 31892 41982
rect 32172 41972 32228 42028
rect 31500 41356 31668 41412
rect 31500 40964 31556 40974
rect 31500 40626 31556 40908
rect 31500 40574 31502 40626
rect 31554 40574 31556 40626
rect 31500 40562 31556 40574
rect 31388 40516 31444 40526
rect 31388 40292 31444 40460
rect 31388 40236 31556 40292
rect 31388 40068 31444 40078
rect 31388 39730 31444 40012
rect 31388 39678 31390 39730
rect 31442 39678 31444 39730
rect 31388 39666 31444 39678
rect 31276 39340 31444 39396
rect 30380 39116 30884 39172
rect 31276 39172 31332 39182
rect 30044 39004 30548 39060
rect 30044 38834 30100 39004
rect 30492 38948 30548 39004
rect 30492 38882 30548 38892
rect 31164 38948 31220 38958
rect 30044 38782 30046 38834
rect 30098 38782 30100 38834
rect 30044 38770 30100 38782
rect 30156 38836 30212 38846
rect 30380 38836 30436 38846
rect 30156 38834 30380 38836
rect 30156 38782 30158 38834
rect 30210 38782 30380 38834
rect 30156 38780 30380 38782
rect 30156 38770 30212 38780
rect 30380 38770 30436 38780
rect 30044 38612 30100 38622
rect 30100 38556 30324 38612
rect 30044 38546 30100 38556
rect 30268 38388 30324 38556
rect 29932 38332 30100 38388
rect 29708 38210 29764 38220
rect 29148 38098 29204 38108
rect 29484 38164 29540 38174
rect 29036 37884 29204 37940
rect 28924 37828 28980 37838
rect 28924 37734 28980 37772
rect 28588 37538 28644 37548
rect 28700 37548 28868 37604
rect 29036 37604 29092 37614
rect 28700 37378 28756 37548
rect 28700 37326 28702 37378
rect 28754 37326 28756 37378
rect 28700 37314 28756 37326
rect 28588 37266 28644 37278
rect 28588 37214 28590 37266
rect 28642 37214 28644 37266
rect 28588 37156 28644 37214
rect 28812 37268 28868 37278
rect 29036 37268 29092 37548
rect 28812 37266 29092 37268
rect 28812 37214 28814 37266
rect 28866 37214 29092 37266
rect 28812 37212 29092 37214
rect 28812 37202 28868 37212
rect 28588 37100 28756 37156
rect 28476 36988 28644 37044
rect 28588 36932 28644 36988
rect 28364 36876 28532 36932
rect 28252 36370 28308 36382
rect 28252 36318 28254 36370
rect 28306 36318 28308 36370
rect 28252 36036 28308 36318
rect 28364 36260 28420 36270
rect 28364 36166 28420 36204
rect 28252 35970 28308 35980
rect 28252 35812 28308 35822
rect 28140 35810 28308 35812
rect 28140 35758 28254 35810
rect 28306 35758 28308 35810
rect 28140 35756 28308 35758
rect 27132 35476 27188 35486
rect 26908 34242 26964 34300
rect 26908 34190 26910 34242
rect 26962 34190 26964 34242
rect 26908 34178 26964 34190
rect 27020 34804 27076 34814
rect 26796 33954 26852 33964
rect 26908 33572 26964 33582
rect 26908 33458 26964 33516
rect 26908 33406 26910 33458
rect 26962 33406 26964 33458
rect 26908 33394 26964 33406
rect 26460 33292 26628 33348
rect 26460 33124 26516 33134
rect 26460 33030 26516 33068
rect 26572 32676 26628 33292
rect 27020 32786 27076 34748
rect 27132 34468 27188 35420
rect 27132 34402 27188 34412
rect 27020 32734 27022 32786
rect 27074 32734 27076 32786
rect 27020 32722 27076 32734
rect 27132 33684 27188 33694
rect 26460 32620 26628 32676
rect 26124 31724 26404 31780
rect 25900 31714 25956 31724
rect 26124 31556 26180 31566
rect 25676 31220 25732 31230
rect 25564 31218 25732 31220
rect 25564 31166 25678 31218
rect 25730 31166 25732 31218
rect 25564 31164 25732 31166
rect 25676 31154 25732 31164
rect 26124 31108 26180 31500
rect 26348 31556 26404 31724
rect 26348 31490 26404 31500
rect 26124 31042 26180 31052
rect 26124 30884 26180 30894
rect 26124 30790 26180 30828
rect 25116 30210 25172 30268
rect 25116 30158 25118 30210
rect 25170 30158 25172 30210
rect 25116 30146 25172 30158
rect 24780 29894 24836 29932
rect 23884 29650 24052 29652
rect 23884 29598 23886 29650
rect 23938 29598 24052 29650
rect 23884 29596 24052 29598
rect 23884 29586 23940 29596
rect 26460 27972 26516 32620
rect 26572 32452 26628 32462
rect 26572 32358 26628 32396
rect 27020 31892 27076 31902
rect 27132 31892 27188 33628
rect 27244 32564 27300 35756
rect 27356 35588 27412 35598
rect 27356 35364 27412 35532
rect 27468 35588 27524 35598
rect 27692 35588 27748 35598
rect 27468 35586 27636 35588
rect 27468 35534 27470 35586
rect 27522 35534 27636 35586
rect 27468 35532 27636 35534
rect 27468 35522 27524 35532
rect 27580 35364 27636 35532
rect 27692 35494 27748 35532
rect 27356 35308 27524 35364
rect 27356 35140 27412 35150
rect 27356 32788 27412 35084
rect 27468 34354 27524 35308
rect 28140 35308 28196 35756
rect 28252 35746 28308 35756
rect 27580 35298 27636 35308
rect 27692 35252 27748 35262
rect 27692 34802 27748 35196
rect 28028 35252 28196 35308
rect 28476 35252 28532 36876
rect 28588 36482 28644 36876
rect 28588 36430 28590 36482
rect 28642 36430 28644 36482
rect 28588 36418 28644 36430
rect 28588 35812 28644 35822
rect 28700 35812 28756 37100
rect 28812 36370 28868 36382
rect 29036 36372 29092 37212
rect 28812 36318 28814 36370
rect 28866 36318 28868 36370
rect 28812 36260 28868 36318
rect 28812 36194 28868 36204
rect 28924 36316 29092 36372
rect 28644 35756 28756 35812
rect 28588 35718 28644 35756
rect 28924 35308 28980 36316
rect 29148 36148 29204 37884
rect 29484 37828 29540 38108
rect 29820 38050 29876 38062
rect 29820 37998 29822 38050
rect 29874 37998 29876 38050
rect 29260 37380 29316 37390
rect 29260 37286 29316 37324
rect 27916 35140 27972 35150
rect 28028 35140 28084 35252
rect 28476 35186 28532 35196
rect 28700 35252 28980 35308
rect 29036 36092 29204 36148
rect 29260 36260 29316 36270
rect 27916 35138 28196 35140
rect 27916 35086 27918 35138
rect 27970 35086 28196 35138
rect 27916 35084 28196 35086
rect 27916 35074 27972 35084
rect 27692 34750 27694 34802
rect 27746 34750 27748 34802
rect 27468 34302 27470 34354
rect 27522 34302 27524 34354
rect 27468 34290 27524 34302
rect 27580 34468 27636 34478
rect 27580 34242 27636 34412
rect 27580 34190 27582 34242
rect 27634 34190 27636 34242
rect 27580 34178 27636 34190
rect 27692 33570 27748 34750
rect 27692 33518 27694 33570
rect 27746 33518 27748 33570
rect 27692 33506 27748 33518
rect 27804 34690 27860 34702
rect 27804 34638 27806 34690
rect 27858 34638 27860 34690
rect 27468 33460 27524 33470
rect 27468 33012 27524 33404
rect 27468 32946 27524 32956
rect 27468 32788 27524 32798
rect 27356 32786 27524 32788
rect 27356 32734 27470 32786
rect 27522 32734 27524 32786
rect 27356 32732 27524 32734
rect 27468 32722 27524 32732
rect 27244 32498 27300 32508
rect 27020 31890 27188 31892
rect 27020 31838 27022 31890
rect 27074 31838 27188 31890
rect 27020 31836 27188 31838
rect 27020 31826 27076 31836
rect 26572 31780 26628 31790
rect 26572 31444 26628 31724
rect 26572 31378 26628 31388
rect 26796 31556 26852 31566
rect 26796 31220 26852 31500
rect 26796 31154 26852 31164
rect 27804 29876 27860 34638
rect 27916 34692 27972 34702
rect 27916 34130 27972 34636
rect 28028 34356 28084 34366
rect 28028 34262 28084 34300
rect 27916 34078 27918 34130
rect 27970 34078 27972 34130
rect 27916 34066 27972 34078
rect 28028 33908 28084 33918
rect 27916 33570 27972 33582
rect 27916 33518 27918 33570
rect 27970 33518 27972 33570
rect 27916 33458 27972 33518
rect 27916 33406 27918 33458
rect 27970 33406 27972 33458
rect 27916 33394 27972 33406
rect 27916 32788 27972 32798
rect 28028 32788 28084 33852
rect 28140 33460 28196 35084
rect 28588 34916 28644 34926
rect 28588 34822 28644 34860
rect 28476 34692 28532 34702
rect 28140 33394 28196 33404
rect 28252 34690 28532 34692
rect 28252 34638 28478 34690
rect 28530 34638 28532 34690
rect 28252 34636 28532 34638
rect 27916 32786 28084 32788
rect 27916 32734 27918 32786
rect 27970 32734 28084 32786
rect 27916 32732 28084 32734
rect 27916 32722 27972 32732
rect 28252 30436 28308 34636
rect 28476 34626 28532 34636
rect 28476 34468 28532 34478
rect 28476 34354 28532 34412
rect 28476 34302 28478 34354
rect 28530 34302 28532 34354
rect 28476 34290 28532 34302
rect 28364 33234 28420 33246
rect 28364 33182 28366 33234
rect 28418 33182 28420 33234
rect 28364 33124 28420 33182
rect 28700 33236 28756 35252
rect 28924 34018 28980 34030
rect 28924 33966 28926 34018
rect 28978 33966 28980 34018
rect 28924 33906 28980 33966
rect 28924 33854 28926 33906
rect 28978 33854 28980 33906
rect 28924 33684 28980 33854
rect 29036 33908 29092 36092
rect 29148 35924 29204 35934
rect 29148 35830 29204 35868
rect 29260 35810 29316 36204
rect 29260 35758 29262 35810
rect 29314 35758 29316 35810
rect 29260 35746 29316 35758
rect 29484 35588 29540 37772
rect 29596 37940 29652 37950
rect 29596 37492 29652 37884
rect 29708 37828 29764 37838
rect 29708 37604 29764 37772
rect 29708 37538 29764 37548
rect 29596 37426 29652 37436
rect 29708 37268 29764 37278
rect 29708 37174 29764 37212
rect 29820 37044 29876 37998
rect 30044 38052 30100 38332
rect 30268 38322 30324 38332
rect 30716 38610 30772 38622
rect 30716 38558 30718 38610
rect 30770 38558 30772 38610
rect 30156 38276 30212 38286
rect 30716 38276 30772 38558
rect 31052 38610 31108 38622
rect 31052 38558 31054 38610
rect 31106 38558 31108 38610
rect 31052 38500 31108 38558
rect 31052 38434 31108 38444
rect 30716 38220 31108 38276
rect 30156 38182 30212 38220
rect 30044 37996 30212 38052
rect 30044 37828 30100 37838
rect 30044 37268 30100 37772
rect 30156 37380 30212 37996
rect 30940 38050 30996 38062
rect 30940 37998 30942 38050
rect 30994 37998 30996 38050
rect 30716 37938 30772 37950
rect 30716 37886 30718 37938
rect 30770 37886 30772 37938
rect 30380 37380 30436 37390
rect 30156 37378 30324 37380
rect 30156 37326 30158 37378
rect 30210 37326 30324 37378
rect 30156 37324 30324 37326
rect 30156 37314 30212 37324
rect 30044 37202 30100 37212
rect 29820 36978 29876 36988
rect 29932 37154 29988 37166
rect 29932 37102 29934 37154
rect 29986 37102 29988 37154
rect 29932 36596 29988 37102
rect 29932 36530 29988 36540
rect 30156 36596 30212 36606
rect 29036 33842 29092 33852
rect 29260 35532 29540 35588
rect 29596 36482 29652 36494
rect 29596 36430 29598 36482
rect 29650 36430 29652 36482
rect 29596 35812 29652 36430
rect 29932 36372 29988 36382
rect 30156 36372 30212 36540
rect 29932 36370 30212 36372
rect 29932 36318 29934 36370
rect 29986 36318 30212 36370
rect 29932 36316 30212 36318
rect 29932 36306 29988 36316
rect 29820 36258 29876 36270
rect 29820 36206 29822 36258
rect 29874 36206 29876 36258
rect 29820 35812 29876 36206
rect 30268 35924 30324 37324
rect 30380 37286 30436 37324
rect 30380 36708 30436 36746
rect 30380 36642 30436 36652
rect 30716 36708 30772 37886
rect 30828 37828 30884 37838
rect 30828 37734 30884 37772
rect 30940 37492 30996 37998
rect 30380 36484 30436 36494
rect 30380 36390 30436 36428
rect 30604 36148 30660 36158
rect 30268 35868 30436 35924
rect 29820 35756 30324 35812
rect 28924 33618 28980 33628
rect 28812 33460 28868 33470
rect 28812 33366 28868 33404
rect 28700 33170 28756 33180
rect 28476 33124 28532 33134
rect 28364 33068 28476 33124
rect 28364 32900 28420 32910
rect 28364 32786 28420 32844
rect 28364 32734 28366 32786
rect 28418 32734 28420 32786
rect 28364 32722 28420 32734
rect 28476 32340 28532 33068
rect 29260 33012 29316 35532
rect 29484 35364 29540 35374
rect 29484 34692 29540 35308
rect 29596 34916 29652 35756
rect 29708 35586 29764 35598
rect 29708 35534 29710 35586
rect 29762 35534 29764 35586
rect 29708 35476 29764 35534
rect 29708 35410 29764 35420
rect 29820 35588 29876 35598
rect 29596 34860 29764 34916
rect 29596 34692 29652 34702
rect 29484 34690 29652 34692
rect 29484 34638 29598 34690
rect 29650 34638 29652 34690
rect 29484 34636 29652 34638
rect 29596 34626 29652 34636
rect 29372 34132 29428 34142
rect 29372 34038 29428 34076
rect 29484 33684 29540 33694
rect 29484 33458 29540 33628
rect 29484 33406 29486 33458
rect 29538 33406 29540 33458
rect 29484 33394 29540 33406
rect 29260 32946 29316 32956
rect 28476 32274 28532 32284
rect 29708 32228 29764 34860
rect 29820 34354 29876 35532
rect 30156 35586 30212 35598
rect 30156 35534 30158 35586
rect 30210 35534 30212 35586
rect 30156 35364 30212 35534
rect 29932 35140 29988 35150
rect 29932 35026 29988 35084
rect 29932 34974 29934 35026
rect 29986 34974 29988 35026
rect 29932 34962 29988 34974
rect 30156 35138 30212 35308
rect 30156 35086 30158 35138
rect 30210 35086 30212 35138
rect 30156 34804 30212 35086
rect 30044 34748 30212 34804
rect 30044 34580 30100 34748
rect 30268 34692 30324 35756
rect 30380 35474 30436 35868
rect 30604 35922 30660 36092
rect 30604 35870 30606 35922
rect 30658 35870 30660 35922
rect 30604 35858 30660 35870
rect 30716 35700 30772 36652
rect 30828 37436 30996 37492
rect 30828 36596 30884 37436
rect 30940 37266 30996 37278
rect 30940 37214 30942 37266
rect 30994 37214 30996 37266
rect 30940 37156 30996 37214
rect 30940 37090 30996 37100
rect 30884 36540 30996 36596
rect 30828 36530 30884 36540
rect 30380 35422 30382 35474
rect 30434 35422 30436 35474
rect 30380 35410 30436 35422
rect 30604 35644 30772 35700
rect 30828 36258 30884 36270
rect 30828 36206 30830 36258
rect 30882 36206 30884 36258
rect 30492 34916 30548 34926
rect 30492 34822 30548 34860
rect 29820 34302 29822 34354
rect 29874 34302 29876 34354
rect 29820 34244 29876 34302
rect 29820 34178 29876 34188
rect 29932 34524 30100 34580
rect 30156 34636 30324 34692
rect 29708 32162 29764 32172
rect 28252 30370 28308 30380
rect 27804 29810 27860 29820
rect 26460 27906 26516 27916
rect 28588 28196 28644 28206
rect 28588 26404 28644 28140
rect 28588 26338 28644 26348
rect 29932 26292 29988 34524
rect 30156 34468 30212 34636
rect 30044 34412 30212 34468
rect 30380 34580 30436 34590
rect 30044 27524 30100 34412
rect 30380 34354 30436 34524
rect 30380 34302 30382 34354
rect 30434 34302 30436 34354
rect 30380 34290 30436 34302
rect 30156 34244 30212 34254
rect 30156 33906 30212 34188
rect 30156 33854 30158 33906
rect 30210 33854 30212 33906
rect 30156 33842 30212 33854
rect 30044 27458 30100 27468
rect 30268 31668 30324 31678
rect 29932 26226 29988 26236
rect 30268 24724 30324 31612
rect 30604 29540 30660 35644
rect 30828 35364 30884 36206
rect 30828 35298 30884 35308
rect 30940 35252 30996 36540
rect 30940 35186 30996 35196
rect 30940 35028 30996 35038
rect 30940 34934 30996 34972
rect 30716 34356 30772 34366
rect 30716 34262 30772 34300
rect 31052 32788 31108 38220
rect 31164 37492 31220 38892
rect 31276 38946 31332 39116
rect 31276 38894 31278 38946
rect 31330 38894 31332 38946
rect 31276 38882 31332 38894
rect 31276 38500 31332 38510
rect 31276 38276 31332 38444
rect 31276 38210 31332 38220
rect 31276 37938 31332 37950
rect 31276 37886 31278 37938
rect 31330 37886 31332 37938
rect 31276 37828 31332 37886
rect 31276 37762 31332 37772
rect 31276 37492 31332 37502
rect 31164 37490 31332 37492
rect 31164 37438 31278 37490
rect 31330 37438 31332 37490
rect 31164 37436 31332 37438
rect 31276 37426 31332 37436
rect 31388 36706 31444 39340
rect 31500 38052 31556 40236
rect 31500 37986 31556 37996
rect 31388 36654 31390 36706
rect 31442 36654 31444 36706
rect 31388 36594 31444 36654
rect 31388 36542 31390 36594
rect 31442 36542 31444 36594
rect 31388 36530 31444 36542
rect 31500 37492 31556 37502
rect 31500 36372 31556 37436
rect 31612 36708 31668 41356
rect 31724 41188 31780 41198
rect 31836 41188 31892 41916
rect 32060 41916 32228 41972
rect 32060 41746 32116 41916
rect 32060 41694 32062 41746
rect 32114 41694 32116 41746
rect 32060 41636 32116 41694
rect 32060 41570 32116 41580
rect 32284 41746 32340 41758
rect 32284 41694 32286 41746
rect 32338 41694 32340 41746
rect 31724 41186 31892 41188
rect 31724 41134 31726 41186
rect 31778 41134 31892 41186
rect 31724 41132 31892 41134
rect 31724 41122 31780 41132
rect 32284 40964 32340 41694
rect 32284 40898 32340 40908
rect 32396 41188 32452 43148
rect 32732 42980 32788 43374
rect 33068 43428 33124 43932
rect 33516 43428 33572 43438
rect 33068 43362 33124 43372
rect 33180 43426 33572 43428
rect 33180 43374 33518 43426
rect 33570 43374 33572 43426
rect 33180 43372 33572 43374
rect 32732 42914 32788 42924
rect 32844 42754 32900 42766
rect 32844 42702 32846 42754
rect 32898 42702 32900 42754
rect 32508 42532 32564 42542
rect 32508 42438 32564 42476
rect 32844 42196 32900 42702
rect 33068 42644 33124 42654
rect 33068 42550 33124 42588
rect 32844 42130 32900 42140
rect 32620 41860 32676 41870
rect 32508 41746 32564 41758
rect 32508 41694 32510 41746
rect 32562 41694 32564 41746
rect 32508 41636 32564 41694
rect 32508 41570 32564 41580
rect 32620 41746 32676 41804
rect 32620 41694 32622 41746
rect 32674 41694 32676 41746
rect 32284 40516 32340 40526
rect 32284 40290 32340 40460
rect 32284 40238 32286 40290
rect 32338 40238 32340 40290
rect 32284 40226 32340 40238
rect 31948 40178 32004 40190
rect 31948 40126 31950 40178
rect 32002 40126 32004 40178
rect 31948 39732 32004 40126
rect 32060 40180 32116 40190
rect 32060 40086 32116 40124
rect 31948 39666 32004 39676
rect 31724 39618 31780 39630
rect 31724 39566 31726 39618
rect 31778 39566 31780 39618
rect 31724 39396 31780 39566
rect 31724 39330 31780 39340
rect 32396 39172 32452 41132
rect 32620 40964 32676 41694
rect 33180 41412 33236 43372
rect 33516 43362 33572 43372
rect 33516 43204 33572 43214
rect 33516 42980 33572 43148
rect 33516 42914 33572 42924
rect 33180 41346 33236 41356
rect 33292 42644 33348 42654
rect 33292 41748 33348 42588
rect 33628 41972 33684 45052
rect 33852 46004 33908 46014
rect 33740 44660 33796 44670
rect 33740 43204 33796 44604
rect 33852 43652 33908 45948
rect 34188 45892 34244 45902
rect 34076 45890 34244 45892
rect 34076 45838 34190 45890
rect 34242 45838 34244 45890
rect 34076 45836 34244 45838
rect 33964 44994 34020 45006
rect 33964 44942 33966 44994
rect 34018 44942 34020 44994
rect 33964 44546 34020 44942
rect 33964 44494 33966 44546
rect 34018 44494 34020 44546
rect 33964 44434 34020 44494
rect 33964 44382 33966 44434
rect 34018 44382 34020 44434
rect 33964 44370 34020 44382
rect 33964 43652 34020 43662
rect 33852 43650 34020 43652
rect 33852 43598 33966 43650
rect 34018 43598 34020 43650
rect 33852 43596 34020 43598
rect 33964 43586 34020 43596
rect 33740 42642 33796 43148
rect 34076 43092 34132 45836
rect 34188 45826 34244 45836
rect 34076 43026 34132 43036
rect 34188 43314 34244 43326
rect 34188 43262 34190 43314
rect 34242 43262 34244 43314
rect 33740 42590 33742 42642
rect 33794 42590 33796 42642
rect 33740 42578 33796 42590
rect 33964 42642 34020 42654
rect 33964 42590 33966 42642
rect 34018 42590 34020 42642
rect 33068 41188 33124 41198
rect 33068 41094 33124 41132
rect 33292 41074 33348 41692
rect 33404 41916 33684 41972
rect 33852 42530 33908 42542
rect 33852 42478 33854 42530
rect 33906 42478 33908 42530
rect 33404 41636 33460 41916
rect 33404 41570 33460 41580
rect 33516 41748 33572 41758
rect 33292 41022 33294 41074
rect 33346 41022 33348 41074
rect 33292 41010 33348 41022
rect 33404 41188 33460 41198
rect 33404 41074 33460 41132
rect 33404 41022 33406 41074
rect 33458 41022 33460 41074
rect 33404 41010 33460 41022
rect 33516 41074 33572 41692
rect 33516 41022 33518 41074
rect 33570 41022 33572 41074
rect 32620 40898 32676 40908
rect 33180 40964 33236 40974
rect 33180 40870 33236 40908
rect 33516 40740 33572 41022
rect 33628 41746 33684 41758
rect 33628 41694 33630 41746
rect 33682 41694 33684 41746
rect 33628 40964 33684 41694
rect 33852 41076 33908 42478
rect 33964 42532 34020 42590
rect 33964 42466 34020 42476
rect 34188 41970 34244 43262
rect 34300 42868 34356 47292
rect 34860 45220 34916 45230
rect 34860 45126 34916 45164
rect 34412 44994 34468 45006
rect 34412 44942 34414 44994
rect 34466 44942 34468 44994
rect 34412 43876 34468 44942
rect 34636 44546 34692 44558
rect 34636 44494 34638 44546
rect 34690 44494 34692 44546
rect 34524 44100 34580 44110
rect 34524 44006 34580 44044
rect 34412 43810 34468 43820
rect 34412 43428 34468 43438
rect 34636 43428 34692 44494
rect 34972 44098 35028 44110
rect 34972 44046 34974 44098
rect 35026 44046 35028 44098
rect 34972 43988 35028 44046
rect 34972 43922 35028 43932
rect 34860 43876 34916 43886
rect 34860 43764 34916 43820
rect 34860 43708 35028 43764
rect 34412 43426 34692 43428
rect 34412 43374 34414 43426
rect 34466 43374 34692 43426
rect 34412 43372 34692 43374
rect 34748 43540 34804 43550
rect 34412 43362 34468 43372
rect 34524 42980 34580 43372
rect 34748 43204 34804 43484
rect 34748 43138 34804 43148
rect 34860 43426 34916 43438
rect 34860 43374 34862 43426
rect 34914 43374 34916 43426
rect 34860 43092 34916 43374
rect 34860 43026 34916 43036
rect 34412 42868 34468 42878
rect 34300 42866 34468 42868
rect 34300 42814 34414 42866
rect 34466 42814 34468 42866
rect 34524 42848 34580 42924
rect 34300 42812 34468 42814
rect 34412 42802 34468 42812
rect 34972 42644 35028 43708
rect 34972 42578 35028 42588
rect 34860 42532 34916 42542
rect 34188 41918 34190 41970
rect 34242 41918 34244 41970
rect 33964 41748 34020 41758
rect 33964 41746 34132 41748
rect 33964 41694 33966 41746
rect 34018 41694 34132 41746
rect 33964 41692 34132 41694
rect 33964 41682 34020 41692
rect 33852 41010 33908 41020
rect 33628 40898 33684 40908
rect 33404 40684 33572 40740
rect 33404 40628 33460 40684
rect 33628 40628 33684 40638
rect 33404 40562 33460 40572
rect 33516 40572 33628 40628
rect 32732 40516 32788 40526
rect 32956 40516 33012 40526
rect 32788 40460 32956 40516
rect 32732 40450 32788 40460
rect 32956 40450 33012 40460
rect 32620 40404 32676 40414
rect 32620 40292 32676 40348
rect 33516 40292 33572 40572
rect 33628 40562 33684 40572
rect 33964 40404 34020 40414
rect 33964 40310 34020 40348
rect 32620 40236 33572 40292
rect 32508 40180 32564 40218
rect 32508 40114 32564 40124
rect 32508 39956 32564 39966
rect 32508 39842 32564 39900
rect 32508 39790 32510 39842
rect 32562 39790 32564 39842
rect 32508 39778 32564 39790
rect 32620 39396 32676 40236
rect 33628 40180 33684 40190
rect 33516 40178 33684 40180
rect 33516 40126 33630 40178
rect 33682 40126 33684 40178
rect 33516 40124 33684 40126
rect 33068 40068 33124 40078
rect 32396 39106 32452 39116
rect 32508 39340 32676 39396
rect 32732 39732 32788 39742
rect 32172 38948 32228 38958
rect 32172 38854 32228 38892
rect 31724 38834 31780 38846
rect 31724 38782 31726 38834
rect 31778 38782 31780 38834
rect 31724 38500 31780 38782
rect 32396 38836 32452 38846
rect 31948 38724 32004 38762
rect 32396 38742 32452 38780
rect 31948 38658 32004 38668
rect 32508 38610 32564 39340
rect 32732 39284 32788 39676
rect 33068 39730 33124 40012
rect 33068 39678 33070 39730
rect 33122 39678 33124 39730
rect 33068 39666 33124 39678
rect 33180 39732 33236 39742
rect 32844 39620 32900 39630
rect 32844 39618 33012 39620
rect 32844 39566 32846 39618
rect 32898 39566 33012 39618
rect 32844 39564 33012 39566
rect 32844 39554 32900 39564
rect 32508 38558 32510 38610
rect 32562 38558 32564 38610
rect 32508 38546 32564 38558
rect 32620 39228 32788 39284
rect 32956 39284 33012 39564
rect 32956 39228 33124 39284
rect 31724 38434 31780 38444
rect 31948 38500 32004 38510
rect 31836 38388 31892 38398
rect 31724 37154 31780 37166
rect 31724 37102 31726 37154
rect 31778 37102 31780 37154
rect 31724 36932 31780 37102
rect 31724 36866 31780 36876
rect 31612 36642 31668 36652
rect 31388 36316 31556 36372
rect 31724 36372 31780 36382
rect 31276 36148 31332 36158
rect 31276 35924 31332 36092
rect 31276 35858 31332 35868
rect 31164 35588 31220 35598
rect 31164 35586 31332 35588
rect 31164 35534 31166 35586
rect 31218 35534 31332 35586
rect 31164 35532 31332 35534
rect 31164 35522 31220 35532
rect 31164 35252 31220 35262
rect 31164 34354 31220 35196
rect 31164 34302 31166 34354
rect 31218 34302 31220 34354
rect 31164 33684 31220 34302
rect 31164 33618 31220 33628
rect 31276 33908 31332 35532
rect 31388 35026 31444 36316
rect 31724 36278 31780 36316
rect 31612 36260 31668 36270
rect 31612 35924 31668 36204
rect 31612 35858 31668 35868
rect 31500 35700 31556 35710
rect 31500 35606 31556 35644
rect 31836 35474 31892 38332
rect 31948 37938 32004 38444
rect 32172 38276 32228 38286
rect 32396 38276 32452 38286
rect 32620 38276 32676 39228
rect 32844 39172 32900 39182
rect 32900 39116 33012 39172
rect 32844 39106 32900 39116
rect 32732 39060 32788 39070
rect 32732 38948 32788 39004
rect 32844 38948 32900 38958
rect 32732 38946 32900 38948
rect 32732 38894 32846 38946
rect 32898 38894 32900 38946
rect 32732 38892 32900 38894
rect 32844 38882 32900 38892
rect 32172 38274 32452 38276
rect 32172 38222 32174 38274
rect 32226 38222 32398 38274
rect 32450 38222 32452 38274
rect 32172 38220 32452 38222
rect 32172 38210 32228 38220
rect 32396 38210 32452 38220
rect 32508 38220 32676 38276
rect 32732 38610 32788 38622
rect 32732 38558 32734 38610
rect 32786 38558 32788 38610
rect 31948 37886 31950 37938
rect 32002 37886 32004 37938
rect 31948 36372 32004 37886
rect 31948 36306 32004 36316
rect 32060 37826 32116 37838
rect 32060 37774 32062 37826
rect 32114 37774 32116 37826
rect 31948 35924 32004 35934
rect 31948 35830 32004 35868
rect 31836 35422 31838 35474
rect 31890 35422 31892 35474
rect 31388 34974 31390 35026
rect 31442 34974 31444 35026
rect 31388 34962 31444 34974
rect 31724 35028 31780 35038
rect 31836 35028 31892 35422
rect 31724 35026 31892 35028
rect 31724 34974 31726 35026
rect 31778 34974 31892 35026
rect 31724 34972 31892 34974
rect 31724 34962 31780 34972
rect 31276 33572 31332 33852
rect 31276 33506 31332 33516
rect 31052 32722 31108 32732
rect 31948 33460 32004 33470
rect 30604 29474 30660 29484
rect 30268 24658 30324 24668
rect 31948 18340 32004 33404
rect 32060 24052 32116 37774
rect 32172 37156 32228 37166
rect 32228 37100 32340 37156
rect 32172 37062 32228 37100
rect 32172 36596 32228 36606
rect 32172 36258 32228 36540
rect 32172 36206 32174 36258
rect 32226 36206 32228 36258
rect 32172 36148 32228 36206
rect 32172 36082 32228 36092
rect 32284 34916 32340 37100
rect 32396 35812 32452 35822
rect 32396 35718 32452 35756
rect 32284 34850 32340 34860
rect 32172 34692 32228 34702
rect 32172 34132 32228 34636
rect 32172 34066 32228 34076
rect 32508 31332 32564 38220
rect 32620 38052 32676 38062
rect 32620 37958 32676 37996
rect 32732 37490 32788 38558
rect 32956 38164 33012 39116
rect 33068 38836 33124 39228
rect 33068 38770 33124 38780
rect 33180 38274 33236 39676
rect 33292 39284 33348 39294
rect 33292 39060 33348 39228
rect 33516 39284 33572 40124
rect 33628 40114 33684 40124
rect 33740 39730 33796 39742
rect 33740 39678 33742 39730
rect 33794 39678 33796 39730
rect 33628 39620 33684 39630
rect 33628 39526 33684 39564
rect 33516 39218 33572 39228
rect 33740 39284 33796 39678
rect 33740 39218 33796 39228
rect 33852 39620 33908 39630
rect 33908 39564 34020 39620
rect 33404 39060 33460 39070
rect 33516 39060 33572 39070
rect 33292 39004 33404 39060
rect 33460 39058 33572 39060
rect 33460 39006 33518 39058
rect 33570 39006 33572 39058
rect 33460 39004 33572 39006
rect 33404 38928 33460 39004
rect 33516 38994 33572 39004
rect 33852 38948 33908 39564
rect 33964 39506 34020 39564
rect 33964 39454 33966 39506
rect 34018 39454 34020 39506
rect 33964 39442 34020 39454
rect 33740 38892 33908 38948
rect 33516 38836 33572 38846
rect 33740 38836 33796 38892
rect 33516 38610 33572 38780
rect 33628 38780 33796 38836
rect 33964 38836 34020 38846
rect 33628 38668 33684 38780
rect 33964 38742 34020 38780
rect 33628 38612 33796 38668
rect 33516 38558 33518 38610
rect 33570 38558 33572 38610
rect 33516 38546 33572 38558
rect 33180 38222 33182 38274
rect 33234 38222 33236 38274
rect 33180 38210 33236 38222
rect 33068 38164 33124 38174
rect 32956 38162 33124 38164
rect 32956 38110 33070 38162
rect 33122 38110 33124 38162
rect 32956 38108 33124 38110
rect 33068 38098 33124 38108
rect 33516 37826 33572 37838
rect 33516 37774 33518 37826
rect 33570 37774 33572 37826
rect 33516 37716 33572 37774
rect 33516 37650 33572 37660
rect 33740 37716 33796 38612
rect 34076 38612 34132 41692
rect 34188 41524 34244 41918
rect 34636 42530 34916 42532
rect 34636 42478 34862 42530
rect 34914 42478 34916 42530
rect 34636 42476 34916 42478
rect 34636 41636 34692 42476
rect 34860 42466 34916 42476
rect 34972 42420 35028 42430
rect 34972 42194 35028 42364
rect 34972 42142 34974 42194
rect 35026 42142 35028 42194
rect 34972 42130 35028 42142
rect 34636 41570 34692 41580
rect 34748 42084 34804 42094
rect 34188 41458 34244 41468
rect 34636 41412 34692 41422
rect 34412 41300 34468 41310
rect 34412 41206 34468 41244
rect 34636 41186 34692 41356
rect 34636 41134 34638 41186
rect 34690 41134 34692 41186
rect 34300 40740 34356 40750
rect 34188 40404 34244 40442
rect 34188 40338 34244 40348
rect 34300 39284 34356 40684
rect 34636 40068 34692 41134
rect 34748 40626 34804 42028
rect 34748 40574 34750 40626
rect 34802 40574 34804 40626
rect 34748 40562 34804 40574
rect 34860 42082 34916 42094
rect 34860 42030 34862 42082
rect 34914 42030 34916 42082
rect 34860 41972 34916 42030
rect 35084 41972 35140 49532
rect 35616 49200 35728 49800
rect 37632 49200 37744 49800
rect 38332 49364 38388 49374
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 35644 46002 35700 49200
rect 37324 49028 37380 49038
rect 36988 48804 37044 48814
rect 35644 45950 35646 46002
rect 35698 45950 35700 46002
rect 35644 45938 35700 45950
rect 35868 47796 35924 47806
rect 35644 45556 35700 45566
rect 35308 44996 35364 45006
rect 35308 44994 35588 44996
rect 35308 44942 35310 44994
rect 35362 44942 35588 44994
rect 35308 44940 35588 44942
rect 35308 44930 35364 44940
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35308 44548 35364 44558
rect 35308 44212 35364 44492
rect 35532 44436 35588 44940
rect 35532 44370 35588 44380
rect 35308 44118 35364 44156
rect 35308 43428 35364 43438
rect 35644 43428 35700 45500
rect 35756 44994 35812 45006
rect 35756 44942 35758 44994
rect 35810 44942 35812 44994
rect 35756 44436 35812 44942
rect 35756 44370 35812 44380
rect 35756 44098 35812 44110
rect 35756 44046 35758 44098
rect 35810 44046 35812 44098
rect 35756 43652 35812 44046
rect 35756 43586 35812 43596
rect 35756 43428 35812 43438
rect 35308 43426 35476 43428
rect 35308 43374 35310 43426
rect 35362 43374 35476 43426
rect 35308 43372 35476 43374
rect 35644 43426 35812 43428
rect 35644 43374 35758 43426
rect 35810 43374 35812 43426
rect 35644 43372 35812 43374
rect 35308 43362 35364 43372
rect 35420 43314 35476 43372
rect 35756 43362 35812 43372
rect 35420 43262 35422 43314
rect 35474 43262 35476 43314
rect 35420 43250 35476 43262
rect 35756 43204 35812 43214
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35532 42980 35588 42990
rect 35756 42980 35812 43148
rect 35588 42924 35812 42980
rect 35532 42914 35588 42924
rect 35252 42868 35308 42878
rect 35252 42756 35308 42812
rect 35644 42756 35700 42766
rect 35252 42700 35644 42756
rect 35644 42690 35700 42700
rect 35756 42756 35812 42766
rect 35868 42756 35924 47740
rect 36316 47572 36372 47582
rect 36204 47124 36260 47134
rect 36092 45892 36148 45902
rect 36092 45798 36148 45836
rect 36204 45330 36260 47068
rect 36204 45278 36206 45330
rect 36258 45278 36260 45330
rect 36204 45266 36260 45278
rect 36204 44100 36260 44110
rect 35756 42754 35924 42756
rect 35756 42702 35758 42754
rect 35810 42702 35924 42754
rect 35756 42700 35924 42702
rect 36092 44098 36260 44100
rect 36092 44046 36206 44098
rect 36258 44046 36260 44098
rect 36092 44044 36260 44046
rect 35756 42690 35812 42700
rect 34860 41916 35140 41972
rect 35308 42530 35364 42542
rect 35308 42478 35310 42530
rect 35362 42478 35364 42530
rect 35308 41972 35364 42478
rect 35644 42532 35700 42542
rect 35644 42530 35812 42532
rect 35644 42478 35646 42530
rect 35698 42478 35812 42530
rect 35644 42476 35812 42478
rect 35644 42466 35700 42476
rect 34860 40740 34916 41916
rect 35308 41906 35364 41916
rect 35532 41860 35588 41870
rect 35532 41858 35700 41860
rect 35532 41806 35534 41858
rect 35586 41806 35700 41858
rect 35532 41804 35700 41806
rect 35532 41794 35588 41804
rect 35084 41748 35140 41758
rect 35084 41654 35140 41692
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35644 41524 35700 41804
rect 35644 41458 35700 41468
rect 34972 41298 35028 41310
rect 34972 41246 34974 41298
rect 35026 41246 35028 41298
rect 34972 41188 35028 41246
rect 34972 41122 35028 41132
rect 35196 41300 35252 41310
rect 34636 40002 34692 40012
rect 34300 39218 34356 39228
rect 34412 39956 34468 39966
rect 34412 39058 34468 39900
rect 34860 39842 34916 40684
rect 34860 39790 34862 39842
rect 34914 39790 34916 39842
rect 34860 39778 34916 39790
rect 34972 40964 35028 40974
rect 34636 39506 34692 39518
rect 34636 39454 34638 39506
rect 34690 39454 34692 39506
rect 34412 39006 34414 39058
rect 34466 39006 34468 39058
rect 34412 38994 34468 39006
rect 34524 39394 34580 39406
rect 34524 39342 34526 39394
rect 34578 39342 34580 39394
rect 34076 38546 34132 38556
rect 34188 38948 34244 38958
rect 34188 38610 34244 38892
rect 34188 38558 34190 38610
rect 34242 38558 34244 38610
rect 34188 38546 34244 38558
rect 34524 38388 34580 39342
rect 34524 38322 34580 38332
rect 34076 38274 34132 38286
rect 34076 38222 34078 38274
rect 34130 38222 34132 38274
rect 33964 37940 34020 37950
rect 33964 37846 34020 37884
rect 33740 37650 33796 37660
rect 32732 37438 32734 37490
rect 32786 37438 32788 37490
rect 32732 37426 32788 37438
rect 33964 37380 34020 37390
rect 33964 37286 34020 37324
rect 33516 37268 33572 37278
rect 33516 37174 33572 37212
rect 32956 37044 33012 37054
rect 32508 31266 32564 31276
rect 32620 36932 32676 36942
rect 32620 28756 32676 36876
rect 32732 36820 32788 36830
rect 32732 36594 32788 36764
rect 32732 36542 32734 36594
rect 32786 36542 32788 36594
rect 32732 36530 32788 36542
rect 32844 36260 32900 36270
rect 32732 36148 32788 36158
rect 32732 35700 32788 36092
rect 32844 35922 32900 36204
rect 32844 35870 32846 35922
rect 32898 35870 32900 35922
rect 32844 35858 32900 35870
rect 32732 35644 32900 35700
rect 32732 35252 32788 35262
rect 32732 35138 32788 35196
rect 32732 35086 32734 35138
rect 32786 35086 32788 35138
rect 32732 35074 32788 35086
rect 32732 34690 32788 34702
rect 32732 34638 32734 34690
rect 32786 34638 32788 34690
rect 32732 33460 32788 34638
rect 32732 33394 32788 33404
rect 32844 31780 32900 35644
rect 32844 31714 32900 31724
rect 32620 28690 32676 28700
rect 32956 28084 33012 36988
rect 34076 36594 34132 38222
rect 34636 38052 34692 39454
rect 34412 37828 34468 37838
rect 34076 36542 34078 36594
rect 34130 36542 34132 36594
rect 34076 36530 34132 36542
rect 34300 37826 34468 37828
rect 34300 37774 34414 37826
rect 34466 37774 34468 37826
rect 34300 37772 34468 37774
rect 33516 36372 33572 36382
rect 33068 36258 33124 36270
rect 33068 36206 33070 36258
rect 33122 36206 33124 36258
rect 33068 36036 33124 36206
rect 33068 35970 33124 35980
rect 33516 35922 33572 36316
rect 33516 35870 33518 35922
rect 33570 35870 33572 35922
rect 33516 35858 33572 35870
rect 33628 36258 33684 36270
rect 34300 36260 34356 37772
rect 34412 37762 34468 37772
rect 34524 37380 34580 37390
rect 34412 37156 34468 37166
rect 34412 37062 34468 37100
rect 33628 36206 33630 36258
rect 33682 36206 33684 36258
rect 33628 35700 33684 36206
rect 33628 35634 33684 35644
rect 33852 36204 34356 36260
rect 34412 36258 34468 36270
rect 34412 36206 34414 36258
rect 34466 36206 34468 36258
rect 32956 28018 33012 28028
rect 33852 33348 33908 36204
rect 33852 26852 33908 33292
rect 34412 33012 34468 36206
rect 34412 32946 34468 32956
rect 34524 29764 34580 37324
rect 34636 36706 34692 37996
rect 34636 36654 34638 36706
rect 34690 36654 34692 36706
rect 34636 36642 34692 36654
rect 34748 39396 34804 39406
rect 34748 39172 34804 39340
rect 34748 31220 34804 39116
rect 34860 38722 34916 38734
rect 34860 38670 34862 38722
rect 34914 38670 34916 38722
rect 34860 38164 34916 38670
rect 34972 38668 35028 40908
rect 35196 40740 35252 41244
rect 35756 41300 35812 42476
rect 35980 41858 36036 41870
rect 35980 41806 35982 41858
rect 36034 41806 36036 41858
rect 35980 41746 36036 41806
rect 35980 41694 35982 41746
rect 36034 41694 36036 41746
rect 35980 41682 36036 41694
rect 36092 41300 36148 44044
rect 36204 44034 36260 44044
rect 36204 43426 36260 43438
rect 36204 43374 36206 43426
rect 36258 43374 36260 43426
rect 36204 43092 36260 43374
rect 36204 43026 36260 43036
rect 36204 42868 36260 42878
rect 36316 42868 36372 47516
rect 36988 45332 37044 48748
rect 37100 45668 37156 45678
rect 37100 45574 37156 45612
rect 37212 45444 37268 45454
rect 37100 45332 37156 45342
rect 36988 45330 37156 45332
rect 36988 45278 37102 45330
rect 37154 45278 37156 45330
rect 36988 45276 37156 45278
rect 37100 45266 37156 45276
rect 36652 44996 36708 45006
rect 36652 44994 36820 44996
rect 36652 44942 36654 44994
rect 36706 44942 36820 44994
rect 36652 44940 36820 44942
rect 36652 44930 36708 44940
rect 36652 44100 36708 44110
rect 36652 44006 36708 44044
rect 36652 43426 36708 43438
rect 36652 43374 36654 43426
rect 36706 43374 36708 43426
rect 36652 43316 36708 43374
rect 36652 43250 36708 43260
rect 36204 42866 36372 42868
rect 36204 42814 36206 42866
rect 36258 42814 36372 42866
rect 36204 42812 36372 42814
rect 36204 42802 36260 42812
rect 36652 42756 36708 42766
rect 36652 42662 36708 42700
rect 36764 41972 36820 44940
rect 36988 44882 37044 44894
rect 36988 44830 36990 44882
rect 37042 44830 37044 44882
rect 36876 43876 36932 43886
rect 36876 43204 36932 43820
rect 36876 42194 36932 43148
rect 36876 42142 36878 42194
rect 36930 42142 36932 42194
rect 36876 42130 36932 42142
rect 36764 41906 36820 41916
rect 36428 41860 36484 41870
rect 36428 41858 36596 41860
rect 36428 41806 36430 41858
rect 36482 41806 36596 41858
rect 36428 41804 36596 41806
rect 36428 41794 36484 41804
rect 35756 41244 36036 41300
rect 35532 40964 35588 40974
rect 35532 40870 35588 40908
rect 35196 40674 35252 40684
rect 35420 40852 35476 40862
rect 35420 40628 35476 40796
rect 35644 40852 35700 40862
rect 35532 40628 35588 40638
rect 35420 40626 35588 40628
rect 35420 40574 35534 40626
rect 35586 40574 35588 40626
rect 35420 40572 35588 40574
rect 35532 40562 35588 40572
rect 35084 40402 35140 40414
rect 35084 40350 35086 40402
rect 35138 40350 35140 40402
rect 35084 39844 35140 40350
rect 35644 40404 35700 40796
rect 35644 40338 35700 40348
rect 35756 40180 35812 41244
rect 35532 40124 35812 40180
rect 35868 41074 35924 41086
rect 35868 41022 35870 41074
rect 35922 41022 35924 41074
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35084 39778 35140 39788
rect 35196 39842 35252 39854
rect 35196 39790 35198 39842
rect 35250 39790 35252 39842
rect 35084 39508 35140 39518
rect 35196 39508 35252 39790
rect 35308 39844 35364 39854
rect 35308 39508 35364 39788
rect 35532 39730 35588 40124
rect 35532 39678 35534 39730
rect 35586 39678 35588 39730
rect 35532 39666 35588 39678
rect 35756 39956 35812 39966
rect 35196 39452 35364 39508
rect 35084 39414 35140 39452
rect 35196 39284 35252 39294
rect 35756 39284 35812 39900
rect 35084 39228 35196 39284
rect 35084 38836 35140 39228
rect 35196 39218 35252 39228
rect 35420 39228 35812 39284
rect 35420 39172 35476 39228
rect 35420 39106 35476 39116
rect 35532 39060 35588 39070
rect 35756 39060 35812 39070
rect 35588 39058 35812 39060
rect 35588 39006 35758 39058
rect 35810 39006 35812 39058
rect 35588 39004 35812 39006
rect 35532 38994 35588 39004
rect 35756 38994 35812 39004
rect 35084 38770 35140 38780
rect 35308 38836 35364 38846
rect 35308 38742 35364 38780
rect 35868 38668 35924 41022
rect 35980 40626 36036 41244
rect 36092 41234 36148 41244
rect 36428 40964 36484 40974
rect 36428 40870 36484 40908
rect 35980 40574 35982 40626
rect 36034 40574 36036 40626
rect 35980 40562 36036 40574
rect 36428 40404 36484 40414
rect 36428 40310 36484 40348
rect 34972 38612 35140 38668
rect 34860 38098 34916 38108
rect 34860 37940 34916 37950
rect 34860 37828 34916 37884
rect 34860 37826 35028 37828
rect 34860 37774 34862 37826
rect 34914 37774 35028 37826
rect 34860 37772 35028 37774
rect 34860 37762 34916 37772
rect 34860 37492 34916 37502
rect 34860 37398 34916 37436
rect 34860 36706 34916 36718
rect 34860 36654 34862 36706
rect 34914 36654 34916 36706
rect 34860 36594 34916 36654
rect 34860 36542 34862 36594
rect 34914 36542 34916 36594
rect 34860 36530 34916 36542
rect 34972 34692 35028 37772
rect 34972 34626 35028 34636
rect 34748 31154 34804 31164
rect 34524 29698 34580 29708
rect 35084 29316 35140 38612
rect 35756 38612 35924 38668
rect 35980 39394 36036 39406
rect 35980 39342 35982 39394
rect 36034 39342 36036 39394
rect 35980 38612 36036 39342
rect 36092 39396 36148 39406
rect 36148 39340 36260 39396
rect 36092 39330 36148 39340
rect 36204 39060 36260 39340
rect 36204 38966 36260 39004
rect 36428 39394 36484 39406
rect 36428 39342 36430 39394
rect 36482 39342 36484 39394
rect 36316 38948 36372 38958
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35756 38274 35812 38612
rect 35980 38546 36036 38556
rect 36092 38724 36148 38734
rect 35756 38222 35758 38274
rect 35810 38222 35812 38274
rect 35756 38210 35812 38222
rect 35868 38500 35924 38510
rect 35756 38052 35812 38062
rect 35756 37958 35812 37996
rect 35308 37828 35364 37838
rect 35308 37734 35364 37772
rect 35756 37828 35812 37838
rect 35308 37154 35364 37166
rect 35308 37102 35310 37154
rect 35362 37102 35364 37154
rect 35308 37042 35364 37102
rect 35756 37154 35812 37772
rect 35756 37102 35758 37154
rect 35810 37102 35812 37154
rect 35308 36990 35310 37042
rect 35362 36990 35364 37042
rect 35308 36978 35364 36990
rect 35644 37042 35700 37054
rect 35644 36990 35646 37042
rect 35698 36990 35700 37042
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35644 36148 35700 36990
rect 35644 36082 35700 36092
rect 35196 35308 35460 35318
rect 35756 35308 35812 37102
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35532 35252 35812 35308
rect 35532 34468 35588 35252
rect 35868 34580 35924 38444
rect 36092 38164 36148 38668
rect 36204 38164 36260 38174
rect 36092 38162 36260 38164
rect 36092 38110 36206 38162
rect 36258 38110 36260 38162
rect 36092 38108 36260 38110
rect 36204 38098 36260 38108
rect 35868 34514 35924 34524
rect 35532 34402 35588 34412
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 36316 32788 36372 38892
rect 36428 37604 36484 39342
rect 36428 37538 36484 37548
rect 35644 32732 36372 32788
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35084 29250 35140 29260
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 33852 26786 33908 26796
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 32060 23986 32116 23996
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 31948 18274 32004 18284
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 35644 15092 35700 32732
rect 36092 32564 36148 32574
rect 36092 16772 36148 32508
rect 36540 29652 36596 41804
rect 36764 41746 36820 41758
rect 36764 41694 36766 41746
rect 36818 41694 36820 41746
rect 36652 41188 36708 41198
rect 36652 41094 36708 41132
rect 36652 39172 36708 39182
rect 36652 39058 36708 39116
rect 36652 39006 36654 39058
rect 36706 39006 36708 39058
rect 36652 38994 36708 39006
rect 36652 38274 36708 38286
rect 36652 38222 36654 38274
rect 36706 38222 36708 38274
rect 36652 37826 36708 38222
rect 36652 37774 36654 37826
rect 36706 37774 36708 37826
rect 36652 30996 36708 37774
rect 36652 30930 36708 30940
rect 36764 30884 36820 41694
rect 36876 40290 36932 40302
rect 36876 40238 36878 40290
rect 36930 40238 36932 40290
rect 36876 37268 36932 40238
rect 36876 37202 36932 37212
rect 36988 33124 37044 44830
rect 37100 43764 37156 43774
rect 37212 43764 37268 45388
rect 37100 43762 37268 43764
rect 37100 43710 37102 43762
rect 37154 43710 37268 43762
rect 37100 43708 37268 43710
rect 37100 43698 37156 43708
rect 37324 41970 37380 48972
rect 37436 47684 37492 47694
rect 37436 44434 37492 47628
rect 37548 46452 37604 46462
rect 37548 45220 37604 46396
rect 37660 45780 37716 49200
rect 37884 45780 37940 45790
rect 37660 45778 37940 45780
rect 37660 45726 37886 45778
rect 37938 45726 37940 45778
rect 37660 45724 37940 45726
rect 37884 45714 37940 45724
rect 38332 45332 38388 49308
rect 39648 49200 39760 49800
rect 40992 49200 41104 49800
rect 43008 49200 43120 49800
rect 45024 49200 45136 49800
rect 46368 49200 46480 49800
rect 48384 49200 48496 49800
rect 49728 49200 49840 49800
rect 38444 49140 38500 49150
rect 38444 46002 38500 49084
rect 39228 48580 39284 48590
rect 38444 45950 38446 46002
rect 38498 45950 38500 46002
rect 38444 45938 38500 45950
rect 38892 47908 38948 47918
rect 38892 46002 38948 47852
rect 38892 45950 38894 46002
rect 38946 45950 38948 46002
rect 38892 45938 38948 45950
rect 38444 45332 38500 45342
rect 38332 45330 38500 45332
rect 38332 45278 38446 45330
rect 38498 45278 38500 45330
rect 38332 45276 38500 45278
rect 39228 45332 39284 48524
rect 39452 48244 39508 48254
rect 39340 46452 39396 46462
rect 39340 46002 39396 46396
rect 39340 45950 39342 46002
rect 39394 45950 39396 46002
rect 39340 45938 39396 45950
rect 39340 45332 39396 45342
rect 39228 45330 39396 45332
rect 39228 45278 39342 45330
rect 39394 45278 39396 45330
rect 39228 45276 39396 45278
rect 38444 45266 38500 45276
rect 39340 45266 39396 45276
rect 37548 45164 37716 45220
rect 37548 44996 37604 45006
rect 37548 44902 37604 44940
rect 37436 44382 37438 44434
rect 37490 44382 37492 44434
rect 37436 42756 37492 44382
rect 37548 43426 37604 43438
rect 37548 43374 37550 43426
rect 37602 43374 37604 43426
rect 37548 43316 37604 43374
rect 37548 43250 37604 43260
rect 37436 42700 37604 42756
rect 37324 41918 37326 41970
rect 37378 41918 37380 41970
rect 37324 41906 37380 41918
rect 37436 42530 37492 42542
rect 37436 42478 37438 42530
rect 37490 42478 37492 42530
rect 37436 41860 37492 42478
rect 37436 41794 37492 41804
rect 37436 40964 37492 40974
rect 37436 40870 37492 40908
rect 37548 40404 37604 42700
rect 37660 40628 37716 45164
rect 38220 45108 38276 45118
rect 37996 44994 38052 45006
rect 37996 44942 37998 44994
rect 38050 44942 38052 44994
rect 37772 44884 37828 44894
rect 37772 41970 37828 44828
rect 37996 44882 38052 44942
rect 37996 44830 37998 44882
rect 38050 44830 38052 44882
rect 37996 44818 38052 44830
rect 37884 44098 37940 44110
rect 37884 44046 37886 44098
rect 37938 44046 37940 44098
rect 37884 43876 37940 44046
rect 37884 43810 37940 43820
rect 38108 43764 38164 43774
rect 37996 43540 38052 43550
rect 37996 43446 38052 43484
rect 37996 42868 38052 42878
rect 38108 42868 38164 43708
rect 37996 42866 38164 42868
rect 37996 42814 37998 42866
rect 38050 42814 38164 42866
rect 37996 42812 38164 42814
rect 37996 42802 38052 42812
rect 38108 42532 38164 42812
rect 38108 42466 38164 42476
rect 38220 42194 38276 45052
rect 38892 44996 38948 45006
rect 38892 44994 39172 44996
rect 38892 44942 38894 44994
rect 38946 44942 39172 44994
rect 38892 44940 39172 44942
rect 38892 44930 38948 44940
rect 38332 44884 38388 44894
rect 38332 44434 38388 44828
rect 38332 44382 38334 44434
rect 38386 44382 38388 44434
rect 38332 44370 38388 44382
rect 38780 44324 38836 44334
rect 38780 44230 38836 44268
rect 38332 44212 38388 44222
rect 38332 43764 38388 44156
rect 38332 43698 38388 43708
rect 38668 44212 38724 44222
rect 38668 43708 38724 44156
rect 38892 43764 38948 43802
rect 39116 43708 39172 44940
rect 39452 44436 39508 48188
rect 39564 47572 39620 47582
rect 39564 45332 39620 47516
rect 39676 45780 39732 49200
rect 40684 48356 40740 48366
rect 40348 47124 40404 47134
rect 39900 45780 39956 45790
rect 39676 45778 39956 45780
rect 39676 45726 39902 45778
rect 39954 45726 39956 45778
rect 39676 45724 39956 45726
rect 39900 45714 39956 45724
rect 39788 45332 39844 45342
rect 39564 45330 39844 45332
rect 39564 45278 39790 45330
rect 39842 45278 39844 45330
rect 39564 45276 39844 45278
rect 39788 45266 39844 45276
rect 40236 44994 40292 45006
rect 40236 44942 40238 44994
rect 40290 44942 40292 44994
rect 39676 44436 39732 44446
rect 39452 44434 39732 44436
rect 39452 44382 39678 44434
rect 39730 44382 39732 44434
rect 39452 44380 39732 44382
rect 38668 43652 38836 43708
rect 38892 43698 38948 43708
rect 38444 43428 38500 43438
rect 38444 43426 38612 43428
rect 38444 43374 38446 43426
rect 38498 43374 38612 43426
rect 38444 43372 38612 43374
rect 38444 43362 38500 43372
rect 38220 42142 38222 42194
rect 38274 42142 38276 42194
rect 38220 42130 38276 42142
rect 38444 42530 38500 42542
rect 38444 42478 38446 42530
rect 38498 42478 38500 42530
rect 38444 42084 38500 42478
rect 38444 42018 38500 42028
rect 37772 41918 37774 41970
rect 37826 41918 37828 41970
rect 37772 41906 37828 41918
rect 38332 41076 38388 41086
rect 38332 40982 38388 41020
rect 37884 40964 37940 40974
rect 37884 40740 37940 40908
rect 37884 40674 37940 40684
rect 37772 40628 37828 40638
rect 37660 40626 37828 40628
rect 37660 40574 37774 40626
rect 37826 40574 37828 40626
rect 37660 40572 37828 40574
rect 37772 40562 37828 40572
rect 38220 40628 38276 40638
rect 38220 40534 38276 40572
rect 37548 40348 37828 40404
rect 37324 40292 37380 40302
rect 37324 40290 37716 40292
rect 37324 40238 37326 40290
rect 37378 40238 37716 40290
rect 37324 40236 37716 40238
rect 37324 40226 37380 40236
rect 37100 39956 37156 39966
rect 37100 39058 37156 39900
rect 37100 39006 37102 39058
rect 37154 39006 37156 39058
rect 37100 38994 37156 39006
rect 37436 39394 37492 39406
rect 37436 39342 37438 39394
rect 37490 39342 37492 39394
rect 37324 38500 37380 38510
rect 37436 38500 37492 39342
rect 37548 38948 37604 38958
rect 37548 38854 37604 38892
rect 37380 38444 37492 38500
rect 37324 38434 37380 38444
rect 36988 33058 37044 33068
rect 37660 31892 37716 40236
rect 37772 39508 37828 40348
rect 37884 40292 37940 40302
rect 37884 39730 37940 40236
rect 37884 39678 37886 39730
rect 37938 39678 37940 39730
rect 37884 39666 37940 39678
rect 38332 39620 38388 39630
rect 38332 39526 38388 39564
rect 37772 39452 38052 39508
rect 37996 32564 38052 39452
rect 38556 35140 38612 43372
rect 38668 42532 38724 42542
rect 38668 42308 38724 42476
rect 38780 42532 38836 43652
rect 39004 43652 39172 43708
rect 39228 44098 39284 44110
rect 39228 44046 39230 44098
rect 39282 44046 39284 44098
rect 39228 43652 39284 44046
rect 38780 42530 38948 42532
rect 38780 42478 38782 42530
rect 38834 42478 38948 42530
rect 38780 42476 38948 42478
rect 38780 42466 38836 42476
rect 38668 42252 38836 42308
rect 38668 41858 38724 41870
rect 38668 41806 38670 41858
rect 38722 41806 38724 41858
rect 38668 40516 38724 41806
rect 38780 41298 38836 42252
rect 38892 41746 38948 42476
rect 38892 41694 38894 41746
rect 38946 41694 38948 41746
rect 38892 41682 38948 41694
rect 38780 41246 38782 41298
rect 38834 41246 38836 41298
rect 38780 41234 38836 41246
rect 38668 40450 38724 40460
rect 38668 40292 38724 40302
rect 38668 40198 38724 40236
rect 38780 39620 38836 39630
rect 38780 39526 38836 39564
rect 39004 35588 39060 43652
rect 39228 43586 39284 43596
rect 39676 43540 39732 44380
rect 40124 44100 40180 44110
rect 39676 43474 39732 43484
rect 39900 44098 40180 44100
rect 39900 44046 40126 44098
rect 40178 44046 40180 44098
rect 39900 44044 40180 44046
rect 39900 43876 39956 44044
rect 40124 44034 40180 44044
rect 39340 43428 39396 43438
rect 39228 43426 39396 43428
rect 39228 43374 39342 43426
rect 39394 43374 39396 43426
rect 39228 43372 39396 43374
rect 39228 42532 39284 43372
rect 39340 43362 39396 43372
rect 39788 43428 39844 43438
rect 39788 43334 39844 43372
rect 39228 42438 39284 42476
rect 39340 42868 39396 42878
rect 39116 41860 39172 41870
rect 39116 41766 39172 41804
rect 39228 40964 39284 40974
rect 39228 40870 39284 40908
rect 39116 40404 39172 40414
rect 39116 40310 39172 40348
rect 39340 36596 39396 42812
rect 39676 42532 39732 42542
rect 39676 42530 39844 42532
rect 39676 42478 39678 42530
rect 39730 42478 39844 42530
rect 39676 42476 39844 42478
rect 39676 42466 39732 42476
rect 39564 41860 39620 41870
rect 39452 41858 39620 41860
rect 39452 41806 39566 41858
rect 39618 41806 39620 41858
rect 39452 41804 39620 41806
rect 39452 38612 39508 41804
rect 39564 41794 39620 41804
rect 39676 41746 39732 41758
rect 39676 41694 39678 41746
rect 39730 41694 39732 41746
rect 39676 41298 39732 41694
rect 39676 41246 39678 41298
rect 39730 41246 39732 41298
rect 39676 41234 39732 41246
rect 39452 38546 39508 38556
rect 39564 40404 39620 40414
rect 39788 40404 39844 42476
rect 39564 40402 39844 40404
rect 39564 40350 39566 40402
rect 39618 40350 39844 40402
rect 39564 40348 39844 40350
rect 39564 38052 39620 40348
rect 39564 37986 39620 37996
rect 39340 36530 39396 36540
rect 39004 35522 39060 35532
rect 38556 35074 38612 35084
rect 37996 32498 38052 32508
rect 39900 31948 39956 43820
rect 40236 43708 40292 44942
rect 40124 43652 40292 43708
rect 40124 42868 40180 43652
rect 40124 42802 40180 42812
rect 40236 43426 40292 43438
rect 40236 43374 40238 43426
rect 40290 43374 40292 43426
rect 40124 42644 40180 42654
rect 40124 42550 40180 42588
rect 40012 41858 40068 41870
rect 40012 41806 40014 41858
rect 40066 41806 40068 41858
rect 40012 38836 40068 41806
rect 40124 41076 40180 41086
rect 40124 40982 40180 41020
rect 40012 38770 40068 38780
rect 40236 34020 40292 43374
rect 40236 33954 40292 33964
rect 39900 31892 40068 31948
rect 37660 31826 37716 31836
rect 36764 30818 36820 30828
rect 36540 29586 36596 29596
rect 36092 16706 36148 16716
rect 37212 26852 37268 26862
rect 35644 15026 35700 15036
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 23772 11666 23828 11676
rect 19628 11330 19684 11340
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 36428 3444 36484 3454
rect 36428 3350 36484 3388
rect 36988 3444 37044 3454
rect 19404 3278 19406 3330
rect 19458 3278 19460 3330
rect 19404 3266 19460 3278
rect 21420 3330 21476 3342
rect 23100 3332 23156 3342
rect 26460 3332 26516 3342
rect 21420 3278 21422 3330
rect 21474 3278 21476 3330
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20860 1762 20916 1774
rect 20860 1710 20862 1762
rect 20914 1710 20916 1762
rect 20860 800 20916 1710
rect 21420 1762 21476 3278
rect 21420 1710 21422 1762
rect 21474 1710 21476 1762
rect 21420 1698 21476 1710
rect 22876 3330 23156 3332
rect 22876 3278 23102 3330
rect 23154 3278 23156 3330
rect 22876 3276 23156 3278
rect 22876 800 22932 3276
rect 23100 3266 23156 3276
rect 26236 3330 26516 3332
rect 26236 3278 26462 3330
rect 26514 3278 26516 3330
rect 26236 3276 26516 3278
rect 26236 800 26292 3276
rect 26460 3266 26516 3276
rect 28252 3332 28308 3342
rect 28252 800 28308 3276
rect 29260 3332 29316 3342
rect 31836 3332 31892 3342
rect 35196 3332 35252 3342
rect 29260 3238 29316 3276
rect 31612 3330 31892 3332
rect 31612 3278 31838 3330
rect 31890 3278 31892 3330
rect 31612 3276 31892 3278
rect 31612 800 31668 3276
rect 31836 3266 31892 3276
rect 34972 3330 35252 3332
rect 34972 3278 35198 3330
rect 35250 3278 35252 3330
rect 34972 3276 35252 3278
rect 34972 800 35028 3276
rect 35196 3266 35252 3276
rect 36988 800 37044 3388
rect 37212 3330 37268 26796
rect 40012 19908 40068 31892
rect 40348 21812 40404 47068
rect 40572 45668 40628 45678
rect 40572 43764 40628 45612
rect 40684 45330 40740 48300
rect 41804 45892 41860 45902
rect 41804 45798 41860 45836
rect 41356 45780 41412 45790
rect 43036 45780 43092 49200
rect 43260 45780 43316 45790
rect 43036 45778 43316 45780
rect 43036 45726 43262 45778
rect 43314 45726 43316 45778
rect 43036 45724 43316 45726
rect 41356 45686 41412 45724
rect 43260 45714 43316 45724
rect 48076 45780 48132 45790
rect 48412 45780 48468 49200
rect 48076 45778 48468 45780
rect 48076 45726 48078 45778
rect 48130 45726 48468 45778
rect 48076 45724 48468 45726
rect 48076 45714 48132 45724
rect 40684 45278 40686 45330
rect 40738 45278 40740 45330
rect 40684 45266 40740 45278
rect 40908 45668 40964 45678
rect 40684 43764 40740 43774
rect 40572 43762 40740 43764
rect 40572 43710 40686 43762
rect 40738 43710 40740 43762
rect 40572 43708 40740 43710
rect 40684 43698 40740 43708
rect 40572 42530 40628 42542
rect 40572 42478 40574 42530
rect 40626 42478 40628 42530
rect 40572 42420 40628 42478
rect 40572 42354 40628 42364
rect 40460 41858 40516 41870
rect 40460 41806 40462 41858
rect 40514 41806 40516 41858
rect 40460 41748 40516 41806
rect 40460 41682 40516 41692
rect 40572 41412 40628 41422
rect 40572 41298 40628 41356
rect 40572 41246 40574 41298
rect 40626 41246 40628 41298
rect 40572 41234 40628 41246
rect 40908 39060 40964 45612
rect 47740 45668 47796 45678
rect 47740 43762 47796 45612
rect 47740 43710 47742 43762
rect 47794 43710 47796 43762
rect 47740 43698 47796 43710
rect 48076 43538 48132 43550
rect 48076 43486 48078 43538
rect 48130 43486 48132 43538
rect 47292 43426 47348 43438
rect 47292 43374 47294 43426
rect 47346 43374 47348 43426
rect 47292 43092 47348 43374
rect 47292 43026 47348 43036
rect 48076 43092 48132 43486
rect 48076 43026 48132 43036
rect 41468 41858 41524 41870
rect 41468 41806 41470 41858
rect 41522 41806 41524 41858
rect 41468 40068 41524 41806
rect 41468 40002 41524 40012
rect 42028 41636 42084 41646
rect 40908 38994 40964 39004
rect 40348 21746 40404 21756
rect 40012 19842 40068 19852
rect 42028 18452 42084 41580
rect 48076 40514 48132 40526
rect 48076 40462 48078 40514
rect 48130 40462 48132 40514
rect 48076 39732 48132 40462
rect 48076 39666 48132 39676
rect 48076 37826 48132 37838
rect 48076 37774 48078 37826
rect 48130 37774 48132 37826
rect 48076 37716 48132 37774
rect 48076 37650 48132 37660
rect 48076 36258 48132 36270
rect 48076 36206 48078 36258
rect 48130 36206 48132 36258
rect 48076 35700 48132 36206
rect 48076 35634 48132 35644
rect 48076 34690 48132 34702
rect 48076 34638 48078 34690
rect 48130 34638 48132 34690
rect 48076 34356 48132 34638
rect 48076 34290 48132 34300
rect 42028 18386 42084 18396
rect 47740 33908 47796 33918
rect 47516 4226 47572 4238
rect 47516 4174 47518 4226
rect 47570 4174 47572 4226
rect 37548 3444 37604 3454
rect 37548 3350 37604 3388
rect 47516 3444 47572 4174
rect 47516 3378 47572 3388
rect 38556 3332 38612 3342
rect 37212 3278 37214 3330
rect 37266 3278 37268 3330
rect 37212 3266 37268 3278
rect 38332 3330 38612 3332
rect 38332 3278 38558 3330
rect 38610 3278 38612 3330
rect 38332 3276 38612 3278
rect 38332 800 38388 3276
rect 38556 3266 38612 3276
rect 41020 3330 41076 3342
rect 42588 3332 42644 3342
rect 43932 3332 43988 3342
rect 45948 3332 46004 3342
rect 41020 3278 41022 3330
rect 41074 3278 41076 3330
rect 40348 1874 40404 1886
rect 40348 1822 40350 1874
rect 40402 1822 40404 1874
rect 40348 800 40404 1822
rect 41020 1874 41076 3278
rect 41020 1822 41022 1874
rect 41074 1822 41076 1874
rect 41020 1810 41076 1822
rect 42364 3330 42644 3332
rect 42364 3278 42590 3330
rect 42642 3278 42644 3330
rect 42364 3276 42644 3278
rect 42364 800 42420 3276
rect 42588 3266 42644 3276
rect 43708 3330 43988 3332
rect 43708 3278 43934 3330
rect 43986 3278 43988 3330
rect 43708 3276 43988 3278
rect 43708 800 43764 3276
rect 43932 3266 43988 3276
rect 45724 3330 46004 3332
rect 45724 3278 45950 3330
rect 46002 3278 46004 3330
rect 45724 3276 46004 3278
rect 45724 800 45780 3276
rect 45948 3266 46004 3276
rect 47180 3330 47236 3342
rect 47180 3278 47182 3330
rect 47234 3278 47236 3330
rect 0 200 112 800
rect 1344 200 1456 800
rect 3360 200 3472 800
rect 4704 200 4816 800
rect 6720 200 6832 800
rect 8736 200 8848 800
rect 10080 200 10192 800
rect 12096 200 12208 800
rect 14112 200 14224 800
rect 15456 200 15568 800
rect 17472 200 17584 800
rect 18816 200 18928 800
rect 20832 200 20944 800
rect 22848 200 22960 800
rect 24192 200 24304 800
rect 26208 200 26320 800
rect 28224 200 28336 800
rect 29568 200 29680 800
rect 31584 200 31696 800
rect 33600 200 33712 800
rect 34944 200 35056 800
rect 36960 200 37072 800
rect 38304 200 38416 800
rect 40320 200 40432 800
rect 42336 200 42448 800
rect 43680 200 43792 800
rect 45696 200 45808 800
rect 47180 756 47236 3278
rect 47740 3330 47796 33852
rect 48076 32674 48132 32686
rect 48076 32622 48078 32674
rect 48130 32622 48132 32674
rect 48076 32340 48132 32622
rect 48076 32274 48132 32284
rect 48076 31554 48132 31566
rect 48076 31502 48078 31554
rect 48130 31502 48132 31554
rect 48076 30996 48132 31502
rect 48076 30930 48132 30940
rect 48076 29538 48132 29550
rect 48076 29486 48078 29538
rect 48130 29486 48132 29538
rect 48076 28980 48132 29486
rect 48076 28914 48132 28924
rect 48076 26852 48132 26862
rect 48076 26758 48132 26796
rect 48076 23714 48132 23726
rect 48076 23662 48078 23714
rect 48130 23662 48132 23714
rect 48076 23604 48132 23662
rect 48076 23538 48132 23548
rect 48076 22146 48132 22158
rect 48076 22094 48078 22146
rect 48130 22094 48132 22146
rect 48076 21588 48132 22094
rect 48076 21522 48132 21532
rect 48076 18564 48132 18574
rect 48076 18470 48132 18508
rect 48076 17442 48132 17454
rect 48076 17390 48078 17442
rect 48130 17390 48132 17442
rect 48076 16884 48132 17390
rect 48076 16818 48132 16828
rect 48076 12852 48132 12862
rect 48076 12758 48132 12796
rect 48076 12290 48132 12302
rect 48076 12238 48078 12290
rect 48130 12238 48132 12290
rect 48076 11508 48132 12238
rect 48076 11442 48132 11452
rect 48076 9602 48132 9614
rect 48076 9550 48078 9602
rect 48130 9550 48132 9602
rect 48076 9492 48132 9550
rect 48076 9426 48132 9436
rect 48076 8034 48132 8046
rect 48076 7982 48078 8034
rect 48130 7982 48132 8034
rect 48076 7476 48132 7982
rect 48076 7410 48132 7420
rect 48076 6466 48132 6478
rect 48076 6414 48078 6466
rect 48130 6414 48132 6466
rect 48076 6132 48132 6414
rect 48076 6066 48132 6076
rect 48076 4452 48132 4462
rect 48076 4450 48244 4452
rect 48076 4398 48078 4450
rect 48130 4398 48244 4450
rect 48076 4396 48244 4398
rect 48076 4386 48132 4396
rect 48076 3444 48132 3454
rect 48076 3350 48132 3388
rect 47740 3278 47742 3330
rect 47794 3278 47796 3330
rect 47740 3266 47796 3278
rect 48188 2100 48244 4396
rect 48188 2034 48244 2044
rect 49084 3444 49140 3454
rect 49084 800 49140 3388
rect 47180 690 47236 700
rect 47712 200 47824 800
rect 49056 200 49168 800
<< via2 >>
rect 3276 49868 3332 49924
rect 700 47292 756 47348
rect 1820 47740 1876 47796
rect 3164 49084 3220 49140
rect 2268 48300 2324 48356
rect 2156 47068 2212 47124
rect 1708 45724 1764 45780
rect 1932 44940 1988 44996
rect 1820 42364 1876 42420
rect 2156 43708 2212 43764
rect 2156 41970 2212 41972
rect 2156 41918 2158 41970
rect 2158 41918 2210 41970
rect 2210 41918 2212 41970
rect 2156 41916 2212 41918
rect 2492 47292 2548 47348
rect 2604 45724 2660 45780
rect 2380 42028 2436 42084
rect 2380 41186 2436 41188
rect 2380 41134 2382 41186
rect 2382 41134 2434 41186
rect 2434 41134 2436 41186
rect 2380 41132 2436 41134
rect 1932 40962 1988 40964
rect 1932 40910 1934 40962
rect 1934 40910 1986 40962
rect 1986 40910 1988 40962
rect 1932 40908 1988 40910
rect 1820 38332 1876 38388
rect 1820 36988 1876 37044
rect 1820 34972 1876 35028
rect 1820 32956 1876 33012
rect 1820 29596 1876 29652
rect 1820 28252 1876 28308
rect 1820 26236 1876 26292
rect 1820 24220 1876 24276
rect 2716 43372 2772 43428
rect 2828 42866 2884 42868
rect 2828 42814 2830 42866
rect 2830 42814 2882 42866
rect 2882 42814 2884 42866
rect 2828 42812 2884 42814
rect 2716 42140 2772 42196
rect 2380 40348 2436 40404
rect 2492 39116 2548 39172
rect 2828 41692 2884 41748
rect 2828 39730 2884 39732
rect 2828 39678 2830 39730
rect 2830 39678 2882 39730
rect 2882 39678 2884 39730
rect 2828 39676 2884 39678
rect 12236 49868 12292 49924
rect 3836 47964 3892 48020
rect 3724 44828 3780 44884
rect 6972 49196 7028 49252
rect 8092 49532 8148 49588
rect 5180 48972 5236 49028
rect 4956 48636 5012 48692
rect 4956 47068 5012 47124
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4284 45276 4340 45332
rect 3388 43260 3444 43316
rect 3164 42140 3220 42196
rect 3276 41468 3332 41524
rect 4620 45330 4676 45332
rect 4620 45278 4622 45330
rect 4622 45278 4674 45330
rect 4674 45278 4676 45330
rect 4620 45276 4676 45278
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4172 44434 4228 44436
rect 4172 44382 4174 44434
rect 4174 44382 4226 44434
rect 4226 44382 4228 44434
rect 4172 44380 4228 44382
rect 4620 44322 4676 44324
rect 4620 44270 4622 44322
rect 4622 44270 4674 44322
rect 4674 44270 4676 44322
rect 4620 44268 4676 44270
rect 4284 44156 4340 44212
rect 4172 43538 4228 43540
rect 4172 43486 4174 43538
rect 4174 43486 4226 43538
rect 4226 43486 4228 43538
rect 4172 43484 4228 43486
rect 4060 42924 4116 42980
rect 4172 42754 4228 42756
rect 4172 42702 4174 42754
rect 4174 42702 4226 42754
rect 4226 42702 4228 42754
rect 4172 42700 4228 42702
rect 3724 42530 3780 42532
rect 3724 42478 3726 42530
rect 3726 42478 3778 42530
rect 3778 42478 3780 42530
rect 3724 42476 3780 42478
rect 3612 42028 3668 42084
rect 3500 41858 3556 41860
rect 3500 41806 3502 41858
rect 3502 41806 3554 41858
rect 3554 41806 3556 41858
rect 3500 41804 3556 41806
rect 3052 40514 3108 40516
rect 3052 40462 3054 40514
rect 3054 40462 3106 40514
rect 3106 40462 3108 40514
rect 3052 40460 3108 40462
rect 3948 41244 4004 41300
rect 4060 41356 4116 41412
rect 3500 40626 3556 40628
rect 3500 40574 3502 40626
rect 3502 40574 3554 40626
rect 3554 40574 3556 40626
rect 3500 40572 3556 40574
rect 2940 38220 2996 38276
rect 3612 40236 3668 40292
rect 2716 37324 2772 37380
rect 2604 36092 2660 36148
rect 3612 39730 3668 39732
rect 3612 39678 3614 39730
rect 3614 39678 3666 39730
rect 3666 39678 3668 39730
rect 3612 39676 3668 39678
rect 3276 39618 3332 39620
rect 3276 39566 3278 39618
rect 3278 39566 3330 39618
rect 3330 39566 3332 39618
rect 3276 39564 3332 39566
rect 3948 40684 4004 40740
rect 4060 40348 4116 40404
rect 4620 43260 4676 43316
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4620 42364 4676 42420
rect 5068 48076 5124 48132
rect 5964 48860 6020 48916
rect 5852 46396 5908 46452
rect 6860 47740 6916 47796
rect 5516 44604 5572 44660
rect 4956 44156 5012 44212
rect 4956 43650 5012 43652
rect 4956 43598 4958 43650
rect 4958 43598 5010 43650
rect 5010 43598 5012 43650
rect 4956 43596 5012 43598
rect 4396 41858 4452 41860
rect 4396 41806 4398 41858
rect 4398 41806 4450 41858
rect 4450 41806 4452 41858
rect 4396 41804 4452 41806
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4172 39228 4228 39284
rect 4172 38834 4228 38836
rect 4172 38782 4174 38834
rect 4174 38782 4226 38834
rect 4226 38782 4228 38834
rect 4172 38780 4228 38782
rect 1932 23324 1988 23380
rect 2044 22876 2100 22932
rect 1820 20860 1876 20916
rect 4060 38162 4116 38164
rect 4060 38110 4062 38162
rect 4062 38110 4114 38162
rect 4114 38110 4116 38162
rect 4060 38108 4116 38110
rect 4396 40402 4452 40404
rect 4396 40350 4398 40402
rect 4398 40350 4450 40402
rect 4450 40350 4452 40402
rect 4396 40348 4452 40350
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4508 39730 4564 39732
rect 4508 39678 4510 39730
rect 4510 39678 4562 39730
rect 4562 39678 4564 39730
rect 4508 39676 4564 39678
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4620 38220 4676 38276
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 5852 44210 5908 44212
rect 5852 44158 5854 44210
rect 5854 44158 5906 44210
rect 5906 44158 5908 44210
rect 5852 44156 5908 44158
rect 6076 47628 6132 47684
rect 6524 47068 6580 47124
rect 6300 45052 6356 45108
rect 6300 44044 6356 44100
rect 5516 43260 5572 43316
rect 5068 40796 5124 40852
rect 5068 39676 5124 39732
rect 5068 39058 5124 39060
rect 5068 39006 5070 39058
rect 5070 39006 5122 39058
rect 5122 39006 5124 39058
rect 5068 39004 5124 39006
rect 4956 38108 5012 38164
rect 5068 37938 5124 37940
rect 5068 37886 5070 37938
rect 5070 37886 5122 37938
rect 5122 37886 5124 37938
rect 5068 37884 5124 37886
rect 4844 36652 4900 36708
rect 5180 35980 5236 36036
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 6188 41916 6244 41972
rect 5964 41692 6020 41748
rect 5628 41356 5684 41412
rect 5628 39900 5684 39956
rect 5404 39228 5460 39284
rect 5516 38722 5572 38724
rect 5516 38670 5518 38722
rect 5518 38670 5570 38722
rect 5570 38670 5572 38722
rect 5516 38668 5572 38670
rect 5292 34524 5348 34580
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 5852 39788 5908 39844
rect 5852 39340 5908 39396
rect 5964 41244 6020 41300
rect 5852 39116 5908 39172
rect 5740 38780 5796 38836
rect 6300 43596 6356 43652
rect 6748 45106 6804 45108
rect 6748 45054 6750 45106
rect 6750 45054 6802 45106
rect 6802 45054 6804 45106
rect 6748 45052 6804 45054
rect 6748 44434 6804 44436
rect 6748 44382 6750 44434
rect 6750 44382 6802 44434
rect 6802 44382 6804 44434
rect 6748 44380 6804 44382
rect 6636 43596 6692 43652
rect 6860 43596 6916 43652
rect 7084 47516 7140 47572
rect 7196 46620 7252 46676
rect 7308 45948 7364 46004
rect 7308 44492 7364 44548
rect 7308 43148 7364 43204
rect 7084 42924 7140 42980
rect 6524 42812 6580 42868
rect 6636 41970 6692 41972
rect 6636 41918 6638 41970
rect 6638 41918 6690 41970
rect 6690 41918 6692 41970
rect 6636 41916 6692 41918
rect 6972 42082 7028 42084
rect 6972 42030 6974 42082
rect 6974 42030 7026 42082
rect 7026 42030 7028 42082
rect 6972 42028 7028 42030
rect 6860 41916 6916 41972
rect 6972 41074 7028 41076
rect 6972 41022 6974 41074
rect 6974 41022 7026 41074
rect 7026 41022 7028 41074
rect 6972 41020 7028 41022
rect 6860 40684 6916 40740
rect 6076 40124 6132 40180
rect 6972 40236 7028 40292
rect 6636 40124 6692 40180
rect 7868 45164 7924 45220
rect 7644 43820 7700 43876
rect 7196 40684 7252 40740
rect 6188 39900 6244 39956
rect 6860 39676 6916 39732
rect 6860 39340 6916 39396
rect 6076 39004 6132 39060
rect 6524 39116 6580 39172
rect 6412 38946 6468 38948
rect 6412 38894 6414 38946
rect 6414 38894 6466 38946
rect 6466 38894 6468 38946
rect 6412 38892 6468 38894
rect 6524 38668 6580 38724
rect 5852 38332 5908 38388
rect 5964 37490 6020 37492
rect 5964 37438 5966 37490
rect 5966 37438 6018 37490
rect 6018 37438 6020 37490
rect 5964 37436 6020 37438
rect 6748 37996 6804 38052
rect 5628 36764 5684 36820
rect 5628 35308 5684 35364
rect 6300 36594 6356 36596
rect 6300 36542 6302 36594
rect 6302 36542 6354 36594
rect 6354 36542 6356 36594
rect 6300 36540 6356 36542
rect 5516 29484 5572 29540
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 6860 37266 6916 37268
rect 6860 37214 6862 37266
rect 6862 37214 6914 37266
rect 6914 37214 6916 37266
rect 6860 37212 6916 37214
rect 7980 45052 8036 45108
rect 7532 40908 7588 40964
rect 7420 40684 7476 40740
rect 7420 39394 7476 39396
rect 7420 39342 7422 39394
rect 7422 39342 7474 39394
rect 7474 39342 7476 39394
rect 7420 39340 7476 39342
rect 7308 38722 7364 38724
rect 7308 38670 7310 38722
rect 7310 38670 7362 38722
rect 7362 38670 7364 38722
rect 7308 38668 7364 38670
rect 7420 38220 7476 38276
rect 7868 42140 7924 42196
rect 7756 41916 7812 41972
rect 7868 40908 7924 40964
rect 7756 40684 7812 40740
rect 7756 40124 7812 40180
rect 7644 39564 7700 39620
rect 7868 40012 7924 40068
rect 10668 49644 10724 49700
rect 9324 48300 9380 48356
rect 8540 47964 8596 48020
rect 8428 47740 8484 47796
rect 8764 47740 8820 47796
rect 8540 47180 8596 47236
rect 8316 47068 8372 47124
rect 8428 46844 8484 46900
rect 8316 46732 8372 46788
rect 8204 45666 8260 45668
rect 8204 45614 8206 45666
rect 8206 45614 8258 45666
rect 8258 45614 8260 45666
rect 8204 45612 8260 45614
rect 8540 45612 8596 45668
rect 8428 44098 8484 44100
rect 8428 44046 8430 44098
rect 8430 44046 8482 44098
rect 8482 44046 8484 44098
rect 8428 44044 8484 44046
rect 8204 43650 8260 43652
rect 8204 43598 8206 43650
rect 8206 43598 8258 43650
rect 8258 43598 8260 43650
rect 8204 43596 8260 43598
rect 8204 42642 8260 42644
rect 8204 42590 8206 42642
rect 8206 42590 8258 42642
rect 8258 42590 8260 42642
rect 8204 42588 8260 42590
rect 8652 43426 8708 43428
rect 8652 43374 8654 43426
rect 8654 43374 8706 43426
rect 8706 43374 8708 43426
rect 8652 43372 8708 43374
rect 7644 39340 7700 39396
rect 7308 37884 7364 37940
rect 7196 37826 7252 37828
rect 7196 37774 7198 37826
rect 7198 37774 7250 37826
rect 7250 37774 7252 37826
rect 7196 37772 7252 37774
rect 7532 37938 7588 37940
rect 7532 37886 7534 37938
rect 7534 37886 7586 37938
rect 7586 37886 7588 37938
rect 7532 37884 7588 37886
rect 7868 39228 7924 39284
rect 7756 39058 7812 39060
rect 7756 39006 7758 39058
rect 7758 39006 7810 39058
rect 7810 39006 7812 39058
rect 7756 39004 7812 39006
rect 7756 38668 7812 38724
rect 7196 37154 7252 37156
rect 7196 37102 7198 37154
rect 7198 37102 7250 37154
rect 7250 37102 7252 37154
rect 7196 37100 7252 37102
rect 7756 37996 7812 38052
rect 6412 36428 6468 36484
rect 6748 36258 6804 36260
rect 6748 36206 6750 36258
rect 6750 36206 6802 36258
rect 6802 36206 6804 36258
rect 6748 36204 6804 36206
rect 7084 34972 7140 35028
rect 7308 35586 7364 35588
rect 7308 35534 7310 35586
rect 7310 35534 7362 35586
rect 7362 35534 7364 35586
rect 7308 35532 7364 35534
rect 6300 27804 6356 27860
rect 6636 33516 6692 33572
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 2940 20076 2996 20132
rect 1820 18844 1876 18900
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 3948 18284 4004 18340
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 1820 17554 1876 17556
rect 1820 17502 1822 17554
rect 1822 17502 1874 17554
rect 1874 17502 1876 17554
rect 1820 17500 1876 17502
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 1820 15484 1876 15540
rect 8204 39394 8260 39396
rect 8204 39342 8206 39394
rect 8206 39342 8258 39394
rect 8258 39342 8260 39394
rect 8204 39340 8260 39342
rect 7980 38668 8036 38724
rect 8092 37884 8148 37940
rect 7868 37436 7924 37492
rect 7980 37100 8036 37156
rect 8204 37154 8260 37156
rect 8204 37102 8206 37154
rect 8206 37102 8258 37154
rect 8258 37102 8260 37154
rect 8204 37100 8260 37102
rect 7532 30492 7588 30548
rect 7756 35586 7812 35588
rect 7756 35534 7758 35586
rect 7758 35534 7810 35586
rect 7810 35534 7812 35586
rect 7756 35532 7812 35534
rect 8092 36540 8148 36596
rect 8204 34972 8260 35028
rect 8428 40514 8484 40516
rect 8428 40462 8430 40514
rect 8430 40462 8482 40514
rect 8482 40462 8484 40514
rect 8428 40460 8484 40462
rect 9100 47292 9156 47348
rect 8988 44098 9044 44100
rect 8988 44046 8990 44098
rect 8990 44046 9042 44098
rect 9042 44046 9044 44098
rect 8988 44044 9044 44046
rect 8764 42476 8820 42532
rect 9100 42642 9156 42644
rect 9100 42590 9102 42642
rect 9102 42590 9154 42642
rect 9154 42590 9156 42642
rect 9100 42588 9156 42590
rect 8988 42476 9044 42532
rect 8652 41356 8708 41412
rect 10556 47628 10612 47684
rect 10556 47180 10612 47236
rect 10332 46284 10388 46340
rect 9772 46172 9828 46228
rect 9884 45052 9940 45108
rect 9772 44716 9828 44772
rect 9772 44492 9828 44548
rect 9324 42530 9380 42532
rect 9324 42478 9326 42530
rect 9326 42478 9378 42530
rect 9378 42478 9380 42530
rect 9324 42476 9380 42478
rect 9212 42028 9268 42084
rect 8764 41916 8820 41972
rect 8652 41186 8708 41188
rect 8652 41134 8654 41186
rect 8654 41134 8706 41186
rect 8706 41134 8708 41186
rect 8652 41132 8708 41134
rect 8876 41858 8932 41860
rect 8876 41806 8878 41858
rect 8878 41806 8930 41858
rect 8930 41806 8932 41858
rect 8876 41804 8932 41806
rect 9548 41804 9604 41860
rect 9436 41580 9492 41636
rect 8988 41244 9044 41300
rect 9324 41298 9380 41300
rect 9324 41246 9326 41298
rect 9326 41246 9378 41298
rect 9378 41246 9380 41298
rect 9324 41244 9380 41246
rect 9100 41132 9156 41188
rect 9436 40796 9492 40852
rect 8652 40178 8708 40180
rect 8652 40126 8654 40178
rect 8654 40126 8706 40178
rect 8706 40126 8708 40178
rect 8652 40124 8708 40126
rect 8764 39340 8820 39396
rect 8876 40236 8932 40292
rect 8540 38108 8596 38164
rect 8428 37938 8484 37940
rect 8428 37886 8430 37938
rect 8430 37886 8482 37938
rect 8482 37886 8484 37938
rect 8428 37884 8484 37886
rect 8652 37548 8708 37604
rect 8428 36594 8484 36596
rect 8428 36542 8430 36594
rect 8430 36542 8482 36594
rect 8482 36542 8484 36594
rect 8428 36540 8484 36542
rect 8652 35698 8708 35700
rect 8652 35646 8654 35698
rect 8654 35646 8706 35698
rect 8706 35646 8708 35698
rect 8652 35644 8708 35646
rect 9100 39842 9156 39844
rect 9100 39790 9102 39842
rect 9102 39790 9154 39842
rect 9154 39790 9156 39842
rect 9100 39788 9156 39790
rect 9100 39340 9156 39396
rect 9212 39004 9268 39060
rect 8988 37324 9044 37380
rect 8876 36594 8932 36596
rect 8876 36542 8878 36594
rect 8878 36542 8930 36594
rect 8930 36542 8932 36594
rect 8876 36540 8932 36542
rect 8988 36204 9044 36260
rect 8876 35026 8932 35028
rect 8876 34974 8878 35026
rect 8878 34974 8930 35026
rect 8930 34974 8932 35026
rect 8876 34972 8932 34974
rect 8764 34300 8820 34356
rect 8316 33628 8372 33684
rect 7980 33516 8036 33572
rect 9100 31276 9156 31332
rect 9436 39394 9492 39396
rect 9436 39342 9438 39394
rect 9438 39342 9490 39394
rect 9490 39342 9492 39394
rect 9436 39340 9492 39342
rect 9324 37884 9380 37940
rect 9324 36370 9380 36372
rect 9324 36318 9326 36370
rect 9326 36318 9378 36370
rect 9378 36318 9380 36370
rect 9324 36316 9380 36318
rect 10220 44492 10276 44548
rect 10780 48860 10836 48916
rect 11116 48412 11172 48468
rect 10892 45836 10948 45892
rect 11004 45778 11060 45780
rect 11004 45726 11006 45778
rect 11006 45726 11058 45778
rect 11058 45726 11060 45778
rect 11004 45724 11060 45726
rect 11676 49196 11732 49252
rect 11676 46060 11732 46116
rect 11788 48076 11844 48132
rect 12124 46956 12180 47012
rect 11452 45836 11508 45892
rect 10892 44940 10948 44996
rect 11228 45500 11284 45556
rect 11116 45218 11172 45220
rect 11116 45166 11118 45218
rect 11118 45166 11170 45218
rect 11170 45166 11172 45218
rect 11116 45164 11172 45166
rect 11788 45666 11844 45668
rect 11788 45614 11790 45666
rect 11790 45614 11842 45666
rect 11842 45614 11844 45666
rect 11788 45612 11844 45614
rect 10556 43932 10612 43988
rect 10668 43762 10724 43764
rect 10668 43710 10670 43762
rect 10670 43710 10722 43762
rect 10722 43710 10724 43762
rect 10668 43708 10724 43710
rect 9996 42866 10052 42868
rect 9996 42814 9998 42866
rect 9998 42814 10050 42866
rect 10050 42814 10052 42866
rect 9996 42812 10052 42814
rect 9884 42700 9940 42756
rect 10444 42476 10500 42532
rect 9884 42082 9940 42084
rect 9884 42030 9886 42082
rect 9886 42030 9938 42082
rect 9938 42030 9940 42082
rect 9884 42028 9940 42030
rect 9996 42252 10052 42308
rect 10556 42252 10612 42308
rect 10668 43372 10724 43428
rect 10444 42140 10500 42196
rect 10668 42140 10724 42196
rect 9772 41804 9828 41860
rect 9884 41746 9940 41748
rect 9884 41694 9886 41746
rect 9886 41694 9938 41746
rect 9938 41694 9940 41746
rect 9884 41692 9940 41694
rect 9660 41132 9716 41188
rect 9660 40348 9716 40404
rect 9996 41020 10052 41076
rect 9884 40572 9940 40628
rect 9884 40348 9940 40404
rect 9772 39004 9828 39060
rect 10108 39788 10164 39844
rect 10220 39340 10276 39396
rect 9996 39116 10052 39172
rect 10332 38892 10388 38948
rect 10220 38834 10276 38836
rect 10220 38782 10222 38834
rect 10222 38782 10274 38834
rect 10274 38782 10276 38834
rect 10220 38780 10276 38782
rect 10332 38668 10388 38724
rect 9996 38108 10052 38164
rect 10332 37938 10388 37940
rect 10332 37886 10334 37938
rect 10334 37886 10386 37938
rect 10386 37886 10388 37938
rect 10332 37884 10388 37886
rect 10556 41244 10612 41300
rect 11452 45052 11508 45108
rect 11676 45052 11732 45108
rect 11452 44828 11508 44884
rect 11340 43708 11396 43764
rect 11564 43708 11620 43764
rect 10556 39788 10612 39844
rect 10780 39506 10836 39508
rect 10780 39454 10782 39506
rect 10782 39454 10834 39506
rect 10834 39454 10836 39506
rect 10780 39452 10836 39454
rect 10892 39340 10948 39396
rect 10556 39004 10612 39060
rect 10668 38108 10724 38164
rect 9996 37660 10052 37716
rect 9884 37436 9940 37492
rect 9548 35196 9604 35252
rect 9660 36988 9716 37044
rect 9436 34412 9492 34468
rect 9884 36988 9940 37044
rect 10108 36764 10164 36820
rect 10220 37436 10276 37492
rect 9772 36316 9828 36372
rect 9772 35756 9828 35812
rect 10220 35586 10276 35588
rect 10220 35534 10222 35586
rect 10222 35534 10274 35586
rect 10274 35534 10276 35586
rect 10220 35532 10276 35534
rect 10556 37042 10612 37044
rect 10556 36990 10558 37042
rect 10558 36990 10610 37042
rect 10610 36990 10612 37042
rect 10556 36988 10612 36990
rect 10780 36988 10836 37044
rect 10444 35980 10500 36036
rect 10780 35922 10836 35924
rect 10780 35870 10782 35922
rect 10782 35870 10834 35922
rect 10834 35870 10836 35922
rect 10780 35868 10836 35870
rect 9884 34636 9940 34692
rect 10332 35084 10388 35140
rect 10668 34690 10724 34692
rect 10668 34638 10670 34690
rect 10670 34638 10722 34690
rect 10722 34638 10724 34690
rect 10668 34636 10724 34638
rect 10556 34018 10612 34020
rect 10556 33966 10558 34018
rect 10558 33966 10610 34018
rect 10610 33966 10612 34018
rect 10556 33964 10612 33966
rect 11228 43538 11284 43540
rect 11228 43486 11230 43538
rect 11230 43486 11282 43538
rect 11282 43486 11284 43538
rect 11228 43484 11284 43486
rect 11452 42588 11508 42644
rect 11340 41468 11396 41524
rect 11340 40124 11396 40180
rect 11116 38444 11172 38500
rect 11004 38332 11060 38388
rect 11340 38332 11396 38388
rect 11452 38444 11508 38500
rect 11228 38220 11284 38276
rect 11788 43932 11844 43988
rect 11676 43484 11732 43540
rect 11788 40012 11844 40068
rect 11116 37884 11172 37940
rect 11340 37884 11396 37940
rect 11676 38444 11732 38500
rect 11004 37212 11060 37268
rect 11004 36652 11060 36708
rect 11228 36370 11284 36372
rect 11228 36318 11230 36370
rect 11230 36318 11282 36370
rect 11282 36318 11284 36370
rect 11228 36316 11284 36318
rect 11116 35644 11172 35700
rect 11004 34748 11060 34804
rect 11004 34412 11060 34468
rect 11004 33740 11060 33796
rect 11228 34914 11284 34916
rect 11228 34862 11230 34914
rect 11230 34862 11282 34914
rect 11282 34862 11284 34914
rect 11228 34860 11284 34862
rect 11116 33516 11172 33572
rect 10892 31724 10948 31780
rect 11788 36988 11844 37044
rect 11676 36204 11732 36260
rect 11788 36092 11844 36148
rect 11676 35586 11732 35588
rect 11676 35534 11678 35586
rect 11678 35534 11730 35586
rect 11730 35534 11732 35586
rect 11676 35532 11732 35534
rect 11564 35084 11620 35140
rect 11564 34524 11620 34580
rect 11340 31612 11396 31668
rect 11676 33458 11732 33460
rect 11676 33406 11678 33458
rect 11678 33406 11730 33458
rect 11730 33406 11732 33458
rect 11676 33404 11732 33406
rect 10668 30604 10724 30660
rect 9212 29708 9268 29764
rect 7756 24108 7812 24164
rect 7308 23212 7364 23268
rect 21532 49868 21588 49924
rect 32060 49868 32116 49924
rect 17948 49532 18004 49588
rect 16828 49308 16884 49364
rect 12236 46396 12292 46452
rect 12348 47180 12404 47236
rect 12684 46844 12740 46900
rect 12348 45612 12404 45668
rect 12460 45388 12516 45444
rect 12348 44882 12404 44884
rect 12348 44830 12350 44882
rect 12350 44830 12402 44882
rect 12402 44830 12404 44882
rect 12348 44828 12404 44830
rect 12124 43932 12180 43988
rect 12348 44604 12404 44660
rect 12572 44044 12628 44100
rect 15708 49084 15764 49140
rect 13804 48972 13860 49028
rect 13468 47964 13524 48020
rect 12796 46284 12852 46340
rect 13356 46396 13412 46452
rect 13356 46172 13412 46228
rect 12908 44994 12964 44996
rect 12908 44942 12910 44994
rect 12910 44942 12962 44994
rect 12962 44942 12964 44994
rect 12908 44940 12964 44942
rect 12908 44322 12964 44324
rect 12908 44270 12910 44322
rect 12910 44270 12962 44322
rect 12962 44270 12964 44322
rect 12908 44268 12964 44270
rect 12348 43708 12404 43764
rect 13244 45276 13300 45332
rect 13580 45890 13636 45892
rect 13580 45838 13582 45890
rect 13582 45838 13634 45890
rect 13634 45838 13636 45890
rect 13580 45836 13636 45838
rect 13468 44828 13524 44884
rect 12012 42812 12068 42868
rect 12684 43036 12740 43092
rect 12124 42140 12180 42196
rect 12124 41468 12180 41524
rect 12236 38444 12292 38500
rect 12348 39788 12404 39844
rect 12460 39452 12516 39508
rect 12796 42252 12852 42308
rect 12572 38444 12628 38500
rect 12684 38668 12740 38724
rect 13132 41692 13188 41748
rect 12908 41244 12964 41300
rect 12908 39788 12964 39844
rect 14588 48748 14644 48804
rect 13916 47458 13972 47460
rect 13916 47406 13918 47458
rect 13918 47406 13970 47458
rect 13970 47406 13972 47458
rect 13916 47404 13972 47406
rect 14140 47404 14196 47460
rect 13804 44210 13860 44212
rect 13804 44158 13806 44210
rect 13806 44158 13858 44210
rect 13858 44158 13860 44210
rect 13804 44156 13860 44158
rect 14028 45106 14084 45108
rect 14028 45054 14030 45106
rect 14030 45054 14082 45106
rect 14082 45054 14084 45106
rect 14028 45052 14084 45054
rect 14028 44604 14084 44660
rect 13692 43596 13748 43652
rect 13468 41692 13524 41748
rect 13468 40796 13524 40852
rect 13468 40572 13524 40628
rect 14028 43538 14084 43540
rect 14028 43486 14030 43538
rect 14030 43486 14082 43538
rect 14082 43486 14084 43538
rect 14028 43484 14084 43486
rect 13692 43260 13748 43316
rect 14364 44716 14420 44772
rect 14364 43036 14420 43092
rect 14476 43484 14532 43540
rect 13916 42364 13972 42420
rect 13580 40460 13636 40516
rect 13804 40962 13860 40964
rect 13804 40910 13806 40962
rect 13806 40910 13858 40962
rect 13858 40910 13860 40962
rect 13804 40908 13860 40910
rect 13580 39506 13636 39508
rect 13580 39454 13582 39506
rect 13582 39454 13634 39506
rect 13634 39454 13636 39506
rect 13580 39452 13636 39454
rect 12908 38892 12964 38948
rect 13020 38780 13076 38836
rect 12684 38556 12740 38612
rect 12572 38050 12628 38052
rect 12572 37998 12574 38050
rect 12574 37998 12626 38050
rect 12626 37998 12628 38050
rect 12572 37996 12628 37998
rect 12236 37548 12292 37604
rect 12236 37324 12292 37380
rect 12348 37212 12404 37268
rect 12012 36876 12068 36932
rect 12012 36258 12068 36260
rect 12012 36206 12014 36258
rect 12014 36206 12066 36258
rect 12066 36206 12068 36258
rect 12012 36204 12068 36206
rect 12012 35420 12068 35476
rect 12124 34524 12180 34580
rect 12124 33458 12180 33460
rect 12124 33406 12126 33458
rect 12126 33406 12178 33458
rect 12178 33406 12180 33458
rect 12124 33404 12180 33406
rect 11900 32732 11956 32788
rect 12348 36204 12404 36260
rect 12572 36764 12628 36820
rect 12572 36428 12628 36484
rect 12572 36092 12628 36148
rect 12460 35756 12516 35812
rect 12684 34860 12740 34916
rect 12572 34690 12628 34692
rect 12572 34638 12574 34690
rect 12574 34638 12626 34690
rect 12626 34638 12628 34690
rect 12572 34636 12628 34638
rect 12460 34354 12516 34356
rect 12460 34302 12462 34354
rect 12462 34302 12514 34354
rect 12514 34302 12516 34354
rect 12460 34300 12516 34302
rect 12460 33852 12516 33908
rect 12572 33628 12628 33684
rect 12348 33292 12404 33348
rect 12236 32620 12292 32676
rect 12572 33180 12628 33236
rect 12236 32450 12292 32452
rect 12236 32398 12238 32450
rect 12238 32398 12290 32450
rect 12290 32398 12292 32450
rect 12236 32396 12292 32398
rect 12572 31948 12628 32004
rect 12908 36204 12964 36260
rect 13020 36092 13076 36148
rect 12908 35980 12964 36036
rect 13356 38722 13412 38724
rect 13356 38670 13358 38722
rect 13358 38670 13410 38722
rect 13410 38670 13412 38722
rect 13356 38668 13412 38670
rect 14812 48748 14868 48804
rect 14812 48412 14868 48468
rect 14700 47628 14756 47684
rect 15260 46620 15316 46676
rect 15260 45388 15316 45444
rect 15148 45276 15204 45332
rect 14588 43596 14644 43652
rect 14588 42028 14644 42084
rect 14700 45164 14756 45220
rect 14140 41244 14196 41300
rect 14028 41074 14084 41076
rect 14028 41022 14030 41074
rect 14030 41022 14082 41074
rect 14082 41022 14084 41074
rect 14028 41020 14084 41022
rect 13916 40236 13972 40292
rect 14476 41298 14532 41300
rect 14476 41246 14478 41298
rect 14478 41246 14530 41298
rect 14530 41246 14532 41298
rect 14476 41244 14532 41246
rect 14588 41186 14644 41188
rect 14588 41134 14590 41186
rect 14590 41134 14642 41186
rect 14642 41134 14644 41186
rect 14588 41132 14644 41134
rect 13916 39564 13972 39620
rect 13804 39228 13860 39284
rect 13916 38780 13972 38836
rect 14028 39004 14084 39060
rect 13692 38220 13748 38276
rect 14476 39564 14532 39620
rect 14812 43650 14868 43652
rect 14812 43598 14814 43650
rect 14814 43598 14866 43650
rect 14866 43598 14868 43650
rect 14812 43596 14868 43598
rect 15036 42812 15092 42868
rect 15372 45052 15428 45108
rect 15372 44268 15428 44324
rect 15148 43708 15204 43764
rect 14812 42364 14868 42420
rect 16828 48972 16884 49028
rect 16492 48636 16548 48692
rect 15708 43932 15764 43988
rect 15596 42028 15652 42084
rect 15148 41244 15204 41300
rect 15260 41356 15316 41412
rect 14812 40402 14868 40404
rect 14812 40350 14814 40402
rect 14814 40350 14866 40402
rect 14866 40350 14868 40402
rect 14812 40348 14868 40350
rect 15820 47852 15876 47908
rect 15820 47180 15876 47236
rect 16044 47234 16100 47236
rect 16044 47182 16046 47234
rect 16046 47182 16098 47234
rect 16098 47182 16100 47234
rect 16044 47180 16100 47182
rect 16044 44156 16100 44212
rect 15820 41356 15876 41412
rect 13692 37938 13748 37940
rect 13692 37886 13694 37938
rect 13694 37886 13746 37938
rect 13746 37886 13748 37938
rect 13692 37884 13748 37886
rect 13804 37548 13860 37604
rect 14364 38444 14420 38500
rect 14028 38108 14084 38164
rect 14140 37884 14196 37940
rect 13468 37100 13524 37156
rect 14028 37324 14084 37380
rect 13244 36204 13300 36260
rect 13356 36764 13412 36820
rect 13132 35980 13188 36036
rect 12796 33740 12852 33796
rect 13020 33292 13076 33348
rect 13020 32956 13076 33012
rect 13244 34130 13300 34132
rect 13244 34078 13246 34130
rect 13246 34078 13298 34130
rect 13298 34078 13300 34130
rect 13244 34076 13300 34078
rect 13804 36540 13860 36596
rect 13804 36204 13860 36260
rect 13692 36092 13748 36148
rect 13468 35644 13524 35700
rect 14028 36482 14084 36484
rect 14028 36430 14030 36482
rect 14030 36430 14082 36482
rect 14082 36430 14084 36482
rect 14028 36428 14084 36430
rect 13468 34412 13524 34468
rect 13804 35196 13860 35252
rect 13804 34802 13860 34804
rect 13804 34750 13806 34802
rect 13806 34750 13858 34802
rect 13858 34750 13860 34802
rect 13804 34748 13860 34750
rect 13692 34412 13748 34468
rect 13580 33404 13636 33460
rect 13356 33292 13412 33348
rect 13580 32844 13636 32900
rect 12348 26236 12404 26292
rect 13804 31388 13860 31444
rect 14252 36876 14308 36932
rect 14588 36540 14644 36596
rect 14476 35922 14532 35924
rect 14476 35870 14478 35922
rect 14478 35870 14530 35922
rect 14530 35870 14532 35922
rect 14476 35868 14532 35870
rect 14364 35420 14420 35476
rect 14700 34802 14756 34804
rect 14700 34750 14702 34802
rect 14702 34750 14754 34802
rect 14754 34750 14756 34802
rect 14700 34748 14756 34750
rect 14812 37548 14868 37604
rect 14252 34300 14308 34356
rect 14028 32450 14084 32452
rect 14028 32398 14030 32450
rect 14030 32398 14082 32450
rect 14082 32398 14084 32450
rect 14028 32396 14084 32398
rect 15036 36092 15092 36148
rect 15036 35698 15092 35700
rect 15036 35646 15038 35698
rect 15038 35646 15090 35698
rect 15090 35646 15092 35698
rect 15036 35644 15092 35646
rect 14924 35196 14980 35252
rect 14924 34300 14980 34356
rect 15260 37212 15316 37268
rect 15372 36652 15428 36708
rect 15708 35868 15764 35924
rect 16940 48412 16996 48468
rect 16940 47740 16996 47796
rect 17836 47740 17892 47796
rect 16940 47516 16996 47572
rect 17388 45948 17444 46004
rect 16492 41132 16548 41188
rect 16604 45836 16660 45892
rect 16604 45388 16660 45444
rect 16156 38220 16212 38276
rect 15596 35698 15652 35700
rect 15596 35646 15598 35698
rect 15598 35646 15650 35698
rect 15650 35646 15652 35698
rect 15596 35644 15652 35646
rect 15596 35308 15652 35364
rect 16044 35644 16100 35700
rect 15820 35084 15876 35140
rect 14924 33964 14980 34020
rect 14700 33628 14756 33684
rect 14588 33234 14644 33236
rect 14588 33182 14590 33234
rect 14590 33182 14642 33234
rect 14642 33182 14644 33234
rect 14588 33180 14644 33182
rect 15036 33346 15092 33348
rect 15036 33294 15038 33346
rect 15038 33294 15090 33346
rect 15090 33294 15092 33346
rect 15036 33292 15092 33294
rect 14924 32786 14980 32788
rect 14924 32734 14926 32786
rect 14926 32734 14978 32786
rect 14978 32734 14980 32786
rect 14924 32732 14980 32734
rect 14476 32284 14532 32340
rect 14700 31554 14756 31556
rect 14700 31502 14702 31554
rect 14702 31502 14754 31554
rect 14754 31502 14756 31554
rect 14700 31500 14756 31502
rect 14140 31164 14196 31220
rect 14812 31218 14868 31220
rect 14812 31166 14814 31218
rect 14814 31166 14866 31218
rect 14866 31166 14868 31218
rect 14812 31164 14868 31166
rect 15036 31164 15092 31220
rect 15932 34636 15988 34692
rect 15820 34524 15876 34580
rect 15932 34188 15988 34244
rect 15484 33458 15540 33460
rect 15484 33406 15486 33458
rect 15486 33406 15538 33458
rect 15538 33406 15540 33458
rect 15484 33404 15540 33406
rect 14812 30716 14868 30772
rect 15148 29932 15204 29988
rect 15820 33516 15876 33572
rect 15372 32562 15428 32564
rect 15372 32510 15374 32562
rect 15374 32510 15426 32562
rect 15426 32510 15428 32562
rect 15372 32508 15428 32510
rect 15260 30044 15316 30100
rect 13916 29820 13972 29876
rect 13132 24892 13188 24948
rect 12908 23660 12964 23716
rect 11676 21756 11732 21812
rect 15820 33068 15876 33124
rect 16492 39788 16548 39844
rect 16716 45052 16772 45108
rect 17724 46002 17780 46004
rect 17724 45950 17726 46002
rect 17726 45950 17778 46002
rect 17778 45950 17780 46002
rect 17724 45948 17780 45950
rect 17052 43484 17108 43540
rect 16940 43260 16996 43316
rect 17052 42588 17108 42644
rect 17276 43372 17332 43428
rect 16716 41804 16772 41860
rect 16940 42028 16996 42084
rect 17052 41468 17108 41524
rect 17388 43148 17444 43204
rect 17388 42866 17444 42868
rect 17388 42814 17390 42866
rect 17390 42814 17442 42866
rect 17442 42814 17444 42866
rect 17388 42812 17444 42814
rect 17724 45106 17780 45108
rect 17724 45054 17726 45106
rect 17726 45054 17778 45106
rect 17778 45054 17780 45106
rect 17724 45052 17780 45054
rect 23212 49308 23268 49364
rect 18060 49084 18116 49140
rect 17612 43372 17668 43428
rect 17724 44268 17780 44324
rect 17948 44322 18004 44324
rect 17948 44270 17950 44322
rect 17950 44270 18002 44322
rect 18002 44270 18004 44322
rect 17948 44268 18004 44270
rect 17836 43596 17892 43652
rect 17948 43372 18004 43428
rect 17836 42028 17892 42084
rect 18172 45724 18228 45780
rect 18284 48972 18340 49028
rect 18956 48636 19012 48692
rect 18060 42140 18116 42196
rect 18508 47292 18564 47348
rect 18396 43650 18452 43652
rect 18396 43598 18398 43650
rect 18398 43598 18450 43650
rect 18450 43598 18452 43650
rect 18396 43596 18452 43598
rect 18172 41916 18228 41972
rect 17276 41020 17332 41076
rect 17388 41244 17444 41300
rect 16716 40796 16772 40852
rect 16492 38108 16548 38164
rect 16604 36988 16660 37044
rect 16604 35922 16660 35924
rect 16604 35870 16606 35922
rect 16606 35870 16658 35922
rect 16658 35870 16660 35922
rect 16604 35868 16660 35870
rect 16268 34748 16324 34804
rect 16604 35474 16660 35476
rect 16604 35422 16606 35474
rect 16606 35422 16658 35474
rect 16658 35422 16660 35474
rect 16604 35420 16660 35422
rect 16156 34524 16212 34580
rect 16492 35138 16548 35140
rect 16492 35086 16494 35138
rect 16494 35086 16546 35138
rect 16546 35086 16548 35138
rect 16492 35084 16548 35086
rect 16380 34524 16436 34580
rect 16828 36540 16884 36596
rect 17052 38332 17108 38388
rect 17500 41186 17556 41188
rect 17500 41134 17502 41186
rect 17502 41134 17554 41186
rect 17554 41134 17556 41186
rect 17500 41132 17556 41134
rect 17612 40684 17668 40740
rect 17388 38162 17444 38164
rect 17388 38110 17390 38162
rect 17390 38110 17442 38162
rect 17442 38110 17444 38162
rect 17388 38108 17444 38110
rect 17276 36540 17332 36596
rect 17388 36764 17444 36820
rect 16940 35698 16996 35700
rect 16940 35646 16942 35698
rect 16942 35646 16994 35698
rect 16994 35646 16996 35698
rect 16940 35644 16996 35646
rect 16716 34412 16772 34468
rect 16716 34130 16772 34132
rect 16716 34078 16718 34130
rect 16718 34078 16770 34130
rect 16770 34078 16772 34130
rect 16716 34076 16772 34078
rect 16604 34018 16660 34020
rect 16604 33966 16606 34018
rect 16606 33966 16658 34018
rect 16658 33966 16660 34018
rect 16604 33964 16660 33966
rect 16268 33068 16324 33124
rect 15596 32620 15652 32676
rect 16156 32956 16212 33012
rect 15708 32060 15764 32116
rect 15596 30994 15652 30996
rect 15596 30942 15598 30994
rect 15598 30942 15650 30994
rect 15650 30942 15652 30994
rect 15596 30940 15652 30942
rect 16156 32172 16212 32228
rect 16044 31666 16100 31668
rect 16044 31614 16046 31666
rect 16046 31614 16098 31666
rect 16098 31614 16100 31666
rect 16044 31612 16100 31614
rect 15820 30604 15876 30660
rect 16380 32956 16436 33012
rect 16268 31948 16324 32004
rect 16044 30156 16100 30212
rect 16380 31778 16436 31780
rect 16380 31726 16382 31778
rect 16382 31726 16434 31778
rect 16434 31726 16436 31778
rect 16380 31724 16436 31726
rect 16380 31276 16436 31332
rect 16716 32956 16772 33012
rect 16828 32786 16884 32788
rect 16828 32734 16830 32786
rect 16830 32734 16882 32786
rect 16882 32734 16884 32786
rect 16828 32732 16884 32734
rect 16716 32674 16772 32676
rect 16716 32622 16718 32674
rect 16718 32622 16770 32674
rect 16770 32622 16772 32674
rect 16716 32620 16772 32622
rect 17052 33740 17108 33796
rect 17052 33292 17108 33348
rect 16828 32284 16884 32340
rect 17052 32284 17108 32340
rect 16716 31836 16772 31892
rect 16604 30604 16660 30660
rect 15484 27468 15540 27524
rect 16604 29260 16660 29316
rect 16940 31388 16996 31444
rect 16940 31164 16996 31220
rect 16828 30604 16884 30660
rect 17388 35196 17444 35252
rect 17612 36764 17668 36820
rect 18172 41020 18228 41076
rect 18732 47068 18788 47124
rect 18620 45218 18676 45220
rect 18620 45166 18622 45218
rect 18622 45166 18674 45218
rect 18674 45166 18676 45218
rect 18620 45164 18676 45166
rect 18844 44940 18900 44996
rect 18844 44044 18900 44100
rect 18396 42140 18452 42196
rect 18732 42028 18788 42084
rect 18396 41970 18452 41972
rect 18396 41918 18398 41970
rect 18398 41918 18450 41970
rect 18450 41918 18452 41970
rect 18396 41916 18452 41918
rect 18060 40402 18116 40404
rect 18060 40350 18062 40402
rect 18062 40350 18114 40402
rect 18114 40350 18116 40402
rect 18060 40348 18116 40350
rect 18284 40402 18340 40404
rect 18284 40350 18286 40402
rect 18286 40350 18338 40402
rect 18338 40350 18340 40402
rect 18284 40348 18340 40350
rect 17836 39564 17892 39620
rect 17724 36204 17780 36260
rect 17500 35420 17556 35476
rect 17388 34972 17444 35028
rect 17388 34524 17444 34580
rect 17276 33516 17332 33572
rect 17276 32620 17332 32676
rect 17388 32732 17444 32788
rect 17388 32508 17444 32564
rect 17836 38108 17892 38164
rect 17724 35810 17780 35812
rect 17724 35758 17726 35810
rect 17726 35758 17778 35810
rect 17778 35758 17780 35810
rect 17724 35756 17780 35758
rect 17724 33740 17780 33796
rect 18060 38108 18116 38164
rect 18060 37884 18116 37940
rect 18060 36988 18116 37044
rect 17948 36594 18004 36596
rect 17948 36542 17950 36594
rect 17950 36542 18002 36594
rect 18002 36542 18004 36594
rect 17948 36540 18004 36542
rect 17948 36316 18004 36372
rect 17948 35756 18004 35812
rect 17948 35474 18004 35476
rect 17948 35422 17950 35474
rect 17950 35422 18002 35474
rect 18002 35422 18004 35474
rect 17948 35420 18004 35422
rect 18284 39676 18340 39732
rect 18172 36092 18228 36148
rect 18284 37996 18340 38052
rect 18172 35756 18228 35812
rect 18060 34300 18116 34356
rect 17612 33122 17668 33124
rect 17612 33070 17614 33122
rect 17614 33070 17666 33122
rect 17666 33070 17668 33122
rect 17612 33068 17668 33070
rect 17500 31500 17556 31556
rect 17276 31164 17332 31220
rect 17724 32450 17780 32452
rect 17724 32398 17726 32450
rect 17726 32398 17778 32450
rect 17778 32398 17780 32450
rect 17724 32396 17780 32398
rect 17724 31948 17780 32004
rect 17836 31836 17892 31892
rect 18060 31836 18116 31892
rect 17836 31276 17892 31332
rect 17164 30940 17220 30996
rect 17948 30940 18004 30996
rect 17724 30882 17780 30884
rect 17724 30830 17726 30882
rect 17726 30830 17778 30882
rect 17778 30830 17780 30882
rect 17724 30828 17780 30830
rect 17164 30380 17220 30436
rect 19852 46732 19908 46788
rect 18956 43820 19012 43876
rect 19516 45276 19572 45332
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 22764 48972 22820 49028
rect 22204 46284 22260 46340
rect 20636 45276 20692 45332
rect 20860 45388 20916 45444
rect 20188 45164 20244 45220
rect 19628 45052 19684 45108
rect 19516 44268 19572 44324
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 20188 43820 20244 43876
rect 19404 43148 19460 43204
rect 18508 40348 18564 40404
rect 18956 42700 19012 42756
rect 18956 42252 19012 42308
rect 18396 37772 18452 37828
rect 18508 38220 18564 38276
rect 18396 37212 18452 37268
rect 18396 36988 18452 37044
rect 18956 40236 19012 40292
rect 19068 42028 19124 42084
rect 18732 39506 18788 39508
rect 18732 39454 18734 39506
rect 18734 39454 18786 39506
rect 18786 39454 18788 39506
rect 18732 39452 18788 39454
rect 18844 39116 18900 39172
rect 18732 37660 18788 37716
rect 18508 35980 18564 36036
rect 18508 35756 18564 35812
rect 18396 35474 18452 35476
rect 18396 35422 18398 35474
rect 18398 35422 18450 35474
rect 18450 35422 18452 35474
rect 18396 35420 18452 35422
rect 18284 34972 18340 35028
rect 18508 34748 18564 34804
rect 18284 34412 18340 34468
rect 18508 33852 18564 33908
rect 18396 33516 18452 33572
rect 18956 37324 19012 37380
rect 18956 36204 19012 36260
rect 19180 41468 19236 41524
rect 19180 40124 19236 40180
rect 19180 39116 19236 39172
rect 19292 39788 19348 39844
rect 18732 33404 18788 33460
rect 19292 36652 19348 36708
rect 18284 31948 18340 32004
rect 18732 33122 18788 33124
rect 18732 33070 18734 33122
rect 18734 33070 18786 33122
rect 18786 33070 18788 33122
rect 18732 33068 18788 33070
rect 20188 42812 20244 42868
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19516 41916 19572 41972
rect 19964 41804 20020 41860
rect 19964 41186 20020 41188
rect 19964 41134 19966 41186
rect 19966 41134 20018 41186
rect 20018 41134 20020 41186
rect 19964 41132 20020 41134
rect 19628 40796 19684 40852
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19628 37996 19684 38052
rect 19852 38668 19908 38724
rect 19516 37436 19572 37492
rect 19404 34188 19460 34244
rect 19516 36428 19572 36484
rect 19292 34076 19348 34132
rect 19404 33628 19460 33684
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 36482 20132 36484
rect 20076 36430 20078 36482
rect 20078 36430 20130 36482
rect 20130 36430 20132 36482
rect 20076 36428 20132 36430
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 20076 35810 20132 35812
rect 20076 35758 20078 35810
rect 20078 35758 20130 35810
rect 20130 35758 20132 35810
rect 20076 35756 20132 35758
rect 20076 34802 20132 34804
rect 20076 34750 20078 34802
rect 20078 34750 20130 34802
rect 20130 34750 20132 34802
rect 20076 34748 20132 34750
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19852 34188 19908 34244
rect 19852 33516 19908 33572
rect 19740 33404 19796 33460
rect 20076 33458 20132 33460
rect 20076 33406 20078 33458
rect 20078 33406 20130 33458
rect 20130 33406 20132 33458
rect 20076 33404 20132 33406
rect 20412 44492 20468 44548
rect 21532 45276 21588 45332
rect 21196 44604 21252 44660
rect 21868 44828 21924 44884
rect 20412 42812 20468 42868
rect 20860 42866 20916 42868
rect 20860 42814 20862 42866
rect 20862 42814 20914 42866
rect 20914 42814 20916 42866
rect 20860 42812 20916 42814
rect 21196 42252 21252 42308
rect 20972 41356 21028 41412
rect 20860 41074 20916 41076
rect 20860 41022 20862 41074
rect 20862 41022 20914 41074
rect 20914 41022 20916 41074
rect 20860 41020 20916 41022
rect 20412 40460 20468 40516
rect 20412 40124 20468 40180
rect 20524 40236 20580 40292
rect 20300 39900 20356 39956
rect 20188 33180 20244 33236
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 18508 32338 18564 32340
rect 18508 32286 18510 32338
rect 18510 32286 18562 32338
rect 18562 32286 18564 32338
rect 18508 32284 18564 32286
rect 18396 31836 18452 31892
rect 18620 31836 18676 31892
rect 18508 31778 18564 31780
rect 18508 31726 18510 31778
rect 18510 31726 18562 31778
rect 18562 31726 18564 31778
rect 18508 31724 18564 31726
rect 18508 31500 18564 31556
rect 18172 30994 18228 30996
rect 18172 30942 18174 30994
rect 18174 30942 18226 30994
rect 18226 30942 18228 30994
rect 18172 30940 18228 30942
rect 18060 30492 18116 30548
rect 17276 30322 17332 30324
rect 17276 30270 17278 30322
rect 17278 30270 17330 30322
rect 17330 30270 17332 30322
rect 17276 30268 17332 30270
rect 17836 30322 17892 30324
rect 17836 30270 17838 30322
rect 17838 30270 17890 30322
rect 17890 30270 17892 30322
rect 17836 30268 17892 30270
rect 19516 32060 19572 32116
rect 19180 31836 19236 31892
rect 18732 31612 18788 31668
rect 19068 31612 19124 31668
rect 19964 31948 20020 32004
rect 20748 40402 20804 40404
rect 20748 40350 20750 40402
rect 20750 40350 20802 40402
rect 20802 40350 20804 40402
rect 20748 40348 20804 40350
rect 20860 39730 20916 39732
rect 20860 39678 20862 39730
rect 20862 39678 20914 39730
rect 20914 39678 20916 39730
rect 20860 39676 20916 39678
rect 20636 39340 20692 39396
rect 21196 41132 21252 41188
rect 21196 40572 21252 40628
rect 21196 39900 21252 39956
rect 21196 39340 21252 39396
rect 20860 38162 20916 38164
rect 20860 38110 20862 38162
rect 20862 38110 20914 38162
rect 20914 38110 20916 38162
rect 20860 38108 20916 38110
rect 20524 36428 20580 36484
rect 20748 37996 20804 38052
rect 20748 36652 20804 36708
rect 21084 35644 21140 35700
rect 20860 33516 20916 33572
rect 20412 32060 20468 32116
rect 20636 33180 20692 33236
rect 20188 31948 20244 32004
rect 19740 31612 19796 31668
rect 19068 31276 19124 31332
rect 19404 31500 19460 31556
rect 19068 31106 19124 31108
rect 19068 31054 19070 31106
rect 19070 31054 19122 31106
rect 19122 31054 19124 31106
rect 19068 31052 19124 31054
rect 19068 30716 19124 30772
rect 19068 30492 19124 30548
rect 18732 29820 18788 29876
rect 18620 29596 18676 29652
rect 19180 30210 19236 30212
rect 19180 30158 19182 30210
rect 19182 30158 19234 30210
rect 19234 30158 19236 30210
rect 19180 30156 19236 30158
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19740 31218 19796 31220
rect 19740 31166 19742 31218
rect 19742 31166 19794 31218
rect 19794 31166 19796 31218
rect 19740 31164 19796 31166
rect 19628 30492 19684 30548
rect 19740 30716 19796 30772
rect 20524 30940 20580 30996
rect 19852 30044 19908 30100
rect 20300 29932 20356 29988
rect 20524 30770 20580 30772
rect 20524 30718 20526 30770
rect 20526 30718 20578 30770
rect 20578 30718 20580 30770
rect 20524 30716 20580 30718
rect 20412 30604 20468 30660
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 16716 26348 16772 26404
rect 18396 24668 18452 24724
rect 19404 29596 19460 29652
rect 19068 23996 19124 24052
rect 16156 16716 16212 16772
rect 15036 16380 15092 16436
rect 6636 15036 6692 15092
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 1820 14140 1876 14196
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 19740 29650 19796 29652
rect 19740 29598 19742 29650
rect 19742 29598 19794 29650
rect 19794 29598 19796 29650
rect 19740 29596 19796 29598
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20524 29820 20580 29876
rect 20860 33068 20916 33124
rect 20748 32172 20804 32228
rect 20748 31948 20804 32004
rect 20972 32172 21028 32228
rect 20972 31500 21028 31556
rect 21084 32060 21140 32116
rect 20748 30492 20804 30548
rect 20860 30380 20916 30436
rect 20748 30268 20804 30324
rect 20860 30156 20916 30212
rect 20860 29820 20916 29876
rect 20972 29708 21028 29764
rect 20860 29596 20916 29652
rect 21644 42700 21700 42756
rect 21420 41692 21476 41748
rect 22204 44380 22260 44436
rect 22428 44716 22484 44772
rect 22540 43932 22596 43988
rect 22204 43596 22260 43652
rect 21980 43036 22036 43092
rect 21420 40572 21476 40628
rect 21532 40348 21588 40404
rect 22092 41970 22148 41972
rect 22092 41918 22094 41970
rect 22094 41918 22146 41970
rect 22146 41918 22148 41970
rect 22092 41916 22148 41918
rect 22652 44828 22708 44884
rect 22092 41692 22148 41748
rect 22316 41916 22372 41972
rect 22204 40460 22260 40516
rect 21644 38556 21700 38612
rect 21644 38050 21700 38052
rect 21644 37998 21646 38050
rect 21646 37998 21698 38050
rect 21698 37998 21700 38050
rect 21644 37996 21700 37998
rect 21980 38556 22036 38612
rect 21868 37884 21924 37940
rect 21644 36594 21700 36596
rect 21644 36542 21646 36594
rect 21646 36542 21698 36594
rect 21698 36542 21700 36594
rect 21644 36540 21700 36542
rect 21308 33516 21364 33572
rect 21308 32732 21364 32788
rect 21756 35084 21812 35140
rect 21644 35026 21700 35028
rect 21644 34974 21646 35026
rect 21646 34974 21698 35026
rect 21698 34974 21700 35026
rect 21644 34972 21700 34974
rect 22092 37772 22148 37828
rect 21980 37660 22036 37716
rect 21980 36764 22036 36820
rect 21980 35084 22036 35140
rect 21980 33740 22036 33796
rect 21868 33180 21924 33236
rect 21196 30940 21252 30996
rect 21308 32396 21364 32452
rect 21532 32338 21588 32340
rect 21532 32286 21534 32338
rect 21534 32286 21586 32338
rect 21586 32286 21588 32338
rect 21532 32284 21588 32286
rect 21532 31388 21588 31444
rect 21644 31836 21700 31892
rect 21308 30044 21364 30100
rect 21196 29820 21252 29876
rect 21084 29484 21140 29540
rect 20860 29260 20916 29316
rect 21980 32508 22036 32564
rect 22204 37548 22260 37604
rect 22652 43596 22708 43652
rect 22652 43148 22708 43204
rect 22988 48802 23044 48804
rect 22988 48750 22990 48802
rect 22990 48750 23042 48802
rect 23042 48750 23044 48802
rect 22988 48748 23044 48750
rect 22316 38556 22372 38612
rect 22652 40236 22708 40292
rect 22876 45948 22932 46004
rect 22988 45218 23044 45220
rect 22988 45166 22990 45218
rect 22990 45166 23042 45218
rect 23042 45166 23044 45218
rect 22988 45164 23044 45166
rect 22876 42028 22932 42084
rect 23100 42028 23156 42084
rect 24892 49644 24948 49700
rect 22764 40012 22820 40068
rect 22428 38108 22484 38164
rect 22316 37100 22372 37156
rect 22428 37938 22484 37940
rect 22428 37886 22430 37938
rect 22430 37886 22482 37938
rect 22482 37886 22484 37938
rect 22428 37884 22484 37886
rect 22764 37660 22820 37716
rect 22428 36988 22484 37044
rect 22540 37324 22596 37380
rect 22428 34972 22484 35028
rect 22204 33516 22260 33572
rect 22316 33404 22372 33460
rect 22988 40236 23044 40292
rect 23100 37042 23156 37044
rect 23100 36990 23102 37042
rect 23102 36990 23154 37042
rect 23154 36990 23156 37042
rect 23100 36988 23156 36990
rect 23324 47404 23380 47460
rect 23660 47292 23716 47348
rect 23884 47292 23940 47348
rect 23660 44044 23716 44100
rect 23548 43372 23604 43428
rect 23772 43036 23828 43092
rect 23324 41804 23380 41860
rect 23548 42476 23604 42532
rect 23436 40684 23492 40740
rect 23324 37996 23380 38052
rect 23884 42028 23940 42084
rect 23660 41132 23716 41188
rect 23436 37772 23492 37828
rect 23100 34130 23156 34132
rect 23100 34078 23102 34130
rect 23102 34078 23154 34130
rect 23154 34078 23156 34130
rect 23100 34076 23156 34078
rect 22876 33852 22932 33908
rect 22988 33740 23044 33796
rect 22204 31554 22260 31556
rect 22204 31502 22206 31554
rect 22206 31502 22258 31554
rect 22258 31502 22260 31554
rect 22204 31500 22260 31502
rect 22540 32674 22596 32676
rect 22540 32622 22542 32674
rect 22542 32622 22594 32674
rect 22594 32622 22596 32674
rect 22540 32620 22596 32622
rect 22652 31948 22708 32004
rect 23212 33404 23268 33460
rect 23548 35196 23604 35252
rect 23548 34748 23604 34804
rect 23548 33906 23604 33908
rect 23548 33854 23550 33906
rect 23550 33854 23602 33906
rect 23602 33854 23604 33906
rect 23548 33852 23604 33854
rect 23436 33740 23492 33796
rect 23884 37548 23940 37604
rect 23772 36594 23828 36596
rect 23772 36542 23774 36594
rect 23774 36542 23826 36594
rect 23826 36542 23828 36594
rect 23772 36540 23828 36542
rect 24220 47068 24276 47124
rect 24108 43538 24164 43540
rect 24108 43486 24110 43538
rect 24110 43486 24162 43538
rect 24162 43486 24164 43538
rect 24108 43484 24164 43486
rect 25788 49756 25844 49812
rect 25788 49420 25844 49476
rect 25564 49026 25620 49028
rect 25564 48974 25566 49026
rect 25566 48974 25618 49026
rect 25618 48974 25620 49026
rect 25564 48972 25620 48974
rect 25788 48972 25844 49028
rect 24892 45164 24948 45220
rect 25676 45724 25732 45780
rect 24556 44434 24612 44436
rect 24556 44382 24558 44434
rect 24558 44382 24610 44434
rect 24610 44382 24612 44434
rect 24556 44380 24612 44382
rect 24556 43538 24612 43540
rect 24556 43486 24558 43538
rect 24558 43486 24610 43538
rect 24610 43486 24612 43538
rect 24556 43484 24612 43486
rect 24444 43372 24500 43428
rect 24556 42754 24612 42756
rect 24556 42702 24558 42754
rect 24558 42702 24610 42754
rect 24610 42702 24612 42754
rect 24556 42700 24612 42702
rect 24220 41244 24276 41300
rect 24444 41916 24500 41972
rect 24780 44716 24836 44772
rect 25004 44716 25060 44772
rect 25340 44380 25396 44436
rect 24556 40684 24612 40740
rect 24444 40348 24500 40404
rect 24108 37996 24164 38052
rect 24556 39564 24612 39620
rect 24444 39452 24500 39508
rect 24556 39116 24612 39172
rect 25116 42700 25172 42756
rect 25340 42924 25396 42980
rect 25116 42140 25172 42196
rect 25228 42476 25284 42532
rect 25116 40348 25172 40404
rect 26124 49756 26180 49812
rect 26012 49532 26068 49588
rect 26236 49532 26292 49588
rect 26012 49084 26068 49140
rect 26572 49196 26628 49252
rect 26460 49026 26516 49028
rect 26460 48974 26462 49026
rect 26462 48974 26514 49026
rect 26514 48974 26516 49026
rect 26460 48972 26516 48974
rect 26012 48748 26068 48804
rect 26572 47964 26628 48020
rect 25900 44434 25956 44436
rect 25900 44382 25902 44434
rect 25902 44382 25954 44434
rect 25954 44382 25956 44434
rect 25900 44380 25956 44382
rect 25788 42364 25844 42420
rect 25788 42140 25844 42196
rect 25228 39900 25284 39956
rect 25340 40124 25396 40180
rect 24892 39452 24948 39508
rect 24444 38668 24500 38724
rect 24220 36876 24276 36932
rect 24668 38892 24724 38948
rect 24892 38722 24948 38724
rect 24892 38670 24894 38722
rect 24894 38670 24946 38722
rect 24946 38670 24948 38722
rect 24892 38668 24948 38670
rect 24444 37100 24500 37156
rect 25004 37884 25060 37940
rect 25116 37548 25172 37604
rect 24556 36652 24612 36708
rect 24668 36988 24724 37044
rect 23884 34972 23940 35028
rect 23772 34802 23828 34804
rect 23772 34750 23774 34802
rect 23774 34750 23826 34802
rect 23826 34750 23828 34802
rect 23772 34748 23828 34750
rect 23884 34524 23940 34580
rect 23996 35308 24052 35364
rect 23660 33740 23716 33796
rect 23772 33570 23828 33572
rect 23772 33518 23774 33570
rect 23774 33518 23826 33570
rect 23826 33518 23828 33570
rect 23772 33516 23828 33518
rect 23660 33404 23716 33460
rect 22876 32620 22932 32676
rect 22988 31836 23044 31892
rect 22652 31778 22708 31780
rect 22652 31726 22654 31778
rect 22654 31726 22706 31778
rect 22706 31726 22708 31778
rect 22652 31724 22708 31726
rect 22428 31612 22484 31668
rect 21644 30716 21700 30772
rect 21980 31276 22036 31332
rect 21644 29314 21700 29316
rect 21644 29262 21646 29314
rect 21646 29262 21698 29314
rect 21698 29262 21700 29314
rect 21644 29260 21700 29262
rect 21532 27804 21588 27860
rect 20412 27356 20468 27412
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 21980 28754 22036 28756
rect 21980 28702 21982 28754
rect 21982 28702 22034 28754
rect 22034 28702 22036 28754
rect 21980 28700 22036 28702
rect 21756 24556 21812 24612
rect 23324 33068 23380 33124
rect 23212 31666 23268 31668
rect 23212 31614 23214 31666
rect 23214 31614 23266 31666
rect 23266 31614 23268 31666
rect 23212 31612 23268 31614
rect 23100 31276 23156 31332
rect 23212 31388 23268 31444
rect 23548 33068 23604 33124
rect 23436 32956 23492 33012
rect 23548 32732 23604 32788
rect 23436 32620 23492 32676
rect 22652 30156 22708 30212
rect 22428 24556 22484 24612
rect 19404 11452 19460 11508
rect 1820 10108 1876 10164
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 9100 9772 9156 9828
rect 1820 8764 1876 8820
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 1820 6748 1876 6804
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 1372 3500 1428 3556
rect 28 2268 84 2324
rect 2156 3554 2212 3556
rect 2156 3502 2158 3554
rect 2158 3502 2210 3554
rect 2210 3502 2212 3554
rect 2156 3500 2212 3502
rect 1820 3388 1876 3444
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 3052 3612 3108 3668
rect 4284 3666 4340 3668
rect 4284 3614 4286 3666
rect 4286 3614 4338 3666
rect 4338 3614 4340 3666
rect 4284 3612 4340 3614
rect 9100 9548 9156 9604
rect 9548 9602 9604 9604
rect 9548 9550 9550 9602
rect 9550 9550 9602 9602
rect 9602 9550 9604 9602
rect 9548 9548 9604 9550
rect 12684 9548 12740 9604
rect 8764 3612 8820 3668
rect 2492 2268 2548 2324
rect 4732 3276 4788 3332
rect 5740 3330 5796 3332
rect 5740 3278 5742 3330
rect 5742 3278 5794 3330
rect 5794 3278 5796 3330
rect 5740 3276 5796 3278
rect 19628 24444 19684 24500
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 22988 30716 23044 30772
rect 23996 33404 24052 33460
rect 23884 33346 23940 33348
rect 23884 33294 23886 33346
rect 23886 33294 23938 33346
rect 23938 33294 23940 33346
rect 23884 33292 23940 33294
rect 23772 33068 23828 33124
rect 24220 35810 24276 35812
rect 24220 35758 24222 35810
rect 24222 35758 24274 35810
rect 24274 35758 24276 35810
rect 24220 35756 24276 35758
rect 24220 34972 24276 35028
rect 24332 35532 24388 35588
rect 24220 34188 24276 34244
rect 24220 33964 24276 34020
rect 24108 33068 24164 33124
rect 24220 33740 24276 33796
rect 23772 32396 23828 32452
rect 23884 32732 23940 32788
rect 23548 31612 23604 31668
rect 23100 29596 23156 29652
rect 22876 29148 22932 29204
rect 22988 28754 23044 28756
rect 22988 28702 22990 28754
rect 22990 28702 23042 28754
rect 23042 28702 23044 28754
rect 22988 28700 23044 28702
rect 23212 28700 23268 28756
rect 22764 26124 22820 26180
rect 22764 19852 22820 19908
rect 22652 18172 22708 18228
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 23436 14812 23492 14868
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 23436 13132 23492 13188
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 23996 32674 24052 32676
rect 23996 32622 23998 32674
rect 23998 32622 24050 32674
rect 24050 32622 24052 32674
rect 23996 32620 24052 32622
rect 24892 35586 24948 35588
rect 24892 35534 24894 35586
rect 24894 35534 24946 35586
rect 24946 35534 24948 35586
rect 24892 35532 24948 35534
rect 25228 37100 25284 37156
rect 25340 37548 25396 37604
rect 25340 36988 25396 37044
rect 25116 34748 25172 34804
rect 24668 34354 24724 34356
rect 24668 34302 24670 34354
rect 24670 34302 24722 34354
rect 24722 34302 24724 34354
rect 24668 34300 24724 34302
rect 25004 34188 25060 34244
rect 24780 34018 24836 34020
rect 24780 33966 24782 34018
rect 24782 33966 24834 34018
rect 24834 33966 24836 34018
rect 24780 33964 24836 33966
rect 24780 33628 24836 33684
rect 25004 33964 25060 34020
rect 24892 33404 24948 33460
rect 25004 33516 25060 33572
rect 24556 33292 24612 33348
rect 24780 33234 24836 33236
rect 24780 33182 24782 33234
rect 24782 33182 24834 33234
rect 24834 33182 24836 33234
rect 24780 33180 24836 33182
rect 24668 32620 24724 32676
rect 24220 32284 24276 32340
rect 24332 32396 24388 32452
rect 23996 31106 24052 31108
rect 23996 31054 23998 31106
rect 23998 31054 24050 31106
rect 24050 31054 24052 31106
rect 23996 31052 24052 31054
rect 23884 30604 23940 30660
rect 23996 30268 24052 30324
rect 23884 30210 23940 30212
rect 23884 30158 23886 30210
rect 23886 30158 23938 30210
rect 23938 30158 23940 30210
rect 23884 30156 23940 30158
rect 24444 30882 24500 30884
rect 24444 30830 24446 30882
rect 24446 30830 24498 30882
rect 24498 30830 24500 30882
rect 24444 30828 24500 30830
rect 24444 30380 24500 30436
rect 24892 32732 24948 32788
rect 25004 32508 25060 32564
rect 25228 36652 25284 36708
rect 25340 36482 25396 36484
rect 25340 36430 25342 36482
rect 25342 36430 25394 36482
rect 25394 36430 25396 36482
rect 25340 36428 25396 36430
rect 25228 35644 25284 35700
rect 25788 40124 25844 40180
rect 25788 38892 25844 38948
rect 25676 38780 25732 38836
rect 25452 35196 25508 35252
rect 25228 34636 25284 34692
rect 25228 32844 25284 32900
rect 25452 34076 25508 34132
rect 25676 35698 25732 35700
rect 25676 35646 25678 35698
rect 25678 35646 25730 35698
rect 25730 35646 25732 35698
rect 25676 35644 25732 35646
rect 25900 38444 25956 38500
rect 25900 37772 25956 37828
rect 25900 37378 25956 37380
rect 25900 37326 25902 37378
rect 25902 37326 25954 37378
rect 25954 37326 25956 37378
rect 25900 37324 25956 37326
rect 26124 42252 26180 42308
rect 27020 48636 27076 48692
rect 30156 48524 30212 48580
rect 28812 48300 28868 48356
rect 27020 47964 27076 48020
rect 27804 47628 27860 47684
rect 27244 47516 27300 47572
rect 26908 45724 26964 45780
rect 27020 46844 27076 46900
rect 27020 45276 27076 45332
rect 26684 44716 26740 44772
rect 26460 41132 26516 41188
rect 26460 40796 26516 40852
rect 26348 38668 26404 38724
rect 26460 40236 26516 40292
rect 26012 37100 26068 37156
rect 26236 38108 26292 38164
rect 26124 36988 26180 37044
rect 26012 36652 26068 36708
rect 26012 36316 26068 36372
rect 25900 36092 25956 36148
rect 25788 34748 25844 34804
rect 25676 34242 25732 34244
rect 25676 34190 25678 34242
rect 25678 34190 25730 34242
rect 25730 34190 25732 34242
rect 25676 34188 25732 34190
rect 25452 33234 25508 33236
rect 25452 33182 25454 33234
rect 25454 33182 25506 33234
rect 25506 33182 25508 33234
rect 25452 33180 25508 33182
rect 25340 31724 25396 31780
rect 25564 32956 25620 33012
rect 25676 32786 25732 32788
rect 25676 32734 25678 32786
rect 25678 32734 25730 32786
rect 25730 32734 25732 32786
rect 25676 32732 25732 32734
rect 25676 31890 25732 31892
rect 25676 31838 25678 31890
rect 25678 31838 25730 31890
rect 25730 31838 25732 31890
rect 25676 31836 25732 31838
rect 26124 35474 26180 35476
rect 26124 35422 26126 35474
rect 26126 35422 26178 35474
rect 26178 35422 26180 35474
rect 26124 35420 26180 35422
rect 26012 34412 26068 34468
rect 26012 33068 26068 33124
rect 26012 32620 26068 32676
rect 25900 31724 25956 31780
rect 26348 36540 26404 36596
rect 26908 41916 26964 41972
rect 26908 41298 26964 41300
rect 26908 41246 26910 41298
rect 26910 41246 26962 41298
rect 26962 41246 26964 41298
rect 26908 41244 26964 41246
rect 27132 45388 27188 45444
rect 26684 39564 26740 39620
rect 27804 47068 27860 47124
rect 27580 46508 27636 46564
rect 27356 45836 27412 45892
rect 27692 46060 27748 46116
rect 28364 46172 28420 46228
rect 28028 46060 28084 46116
rect 27916 45948 27972 46004
rect 27692 45666 27748 45668
rect 27692 45614 27694 45666
rect 27694 45614 27746 45666
rect 27746 45614 27748 45666
rect 27692 45612 27748 45614
rect 27468 45388 27524 45444
rect 27804 45500 27860 45556
rect 27580 44994 27636 44996
rect 27580 44942 27582 44994
rect 27582 44942 27634 44994
rect 27634 44942 27636 44994
rect 27580 44940 27636 44942
rect 27692 43708 27748 43764
rect 27244 39900 27300 39956
rect 27356 41580 27412 41636
rect 27132 39676 27188 39732
rect 26908 38668 26964 38724
rect 26572 35308 26628 35364
rect 26796 36370 26852 36372
rect 26796 36318 26798 36370
rect 26798 36318 26850 36370
rect 26850 36318 26852 36370
rect 26796 36316 26852 36318
rect 27244 39506 27300 39508
rect 27244 39454 27246 39506
rect 27246 39454 27298 39506
rect 27298 39454 27300 39506
rect 27244 39452 27300 39454
rect 27244 39004 27300 39060
rect 27132 37772 27188 37828
rect 27020 37266 27076 37268
rect 27020 37214 27022 37266
rect 27022 37214 27074 37266
rect 27074 37214 27076 37266
rect 27020 37212 27076 37214
rect 27132 36482 27188 36484
rect 27132 36430 27134 36482
rect 27134 36430 27186 36482
rect 27186 36430 27188 36482
rect 27132 36428 27188 36430
rect 27244 36316 27300 36372
rect 27020 35868 27076 35924
rect 28028 45500 28084 45556
rect 28028 45218 28084 45220
rect 28028 45166 28030 45218
rect 28030 45166 28082 45218
rect 28082 45166 28084 45218
rect 28028 45164 28084 45166
rect 28140 45106 28196 45108
rect 28140 45054 28142 45106
rect 28142 45054 28194 45106
rect 28194 45054 28196 45106
rect 28140 45052 28196 45054
rect 28028 44604 28084 44660
rect 27804 43260 27860 43316
rect 27916 42754 27972 42756
rect 27916 42702 27918 42754
rect 27918 42702 27970 42754
rect 27970 42702 27972 42754
rect 27916 42700 27972 42702
rect 27916 41132 27972 41188
rect 28700 45388 28756 45444
rect 28364 44940 28420 44996
rect 29372 48300 29428 48356
rect 28924 47740 28980 47796
rect 29260 45500 29316 45556
rect 29820 47852 29876 47908
rect 29484 47628 29540 47684
rect 28364 44156 28420 44212
rect 28700 44268 28756 44324
rect 28812 44210 28868 44212
rect 28812 44158 28814 44210
rect 28814 44158 28866 44210
rect 28866 44158 28868 44210
rect 28812 44156 28868 44158
rect 28476 42700 28532 42756
rect 29372 44828 29428 44884
rect 29596 45666 29652 45668
rect 29596 45614 29598 45666
rect 29598 45614 29650 45666
rect 29650 45614 29652 45666
rect 29596 45612 29652 45614
rect 30156 47740 30212 47796
rect 30604 48412 30660 48468
rect 30604 47740 30660 47796
rect 30380 47180 30436 47236
rect 30156 45778 30212 45780
rect 30156 45726 30158 45778
rect 30158 45726 30210 45778
rect 30210 45726 30212 45778
rect 30156 45724 30212 45726
rect 29820 45500 29876 45556
rect 30828 48412 30884 48468
rect 30604 46284 30660 46340
rect 30716 47404 30772 47460
rect 30044 45106 30100 45108
rect 30044 45054 30046 45106
rect 30046 45054 30098 45106
rect 30098 45054 30100 45106
rect 30044 45052 30100 45054
rect 29708 44940 29764 44996
rect 30156 44940 30212 44996
rect 29484 44268 29540 44324
rect 29708 44268 29764 44324
rect 29036 43708 29092 43764
rect 29036 43426 29092 43428
rect 29036 43374 29038 43426
rect 29038 43374 29090 43426
rect 29090 43374 29092 43426
rect 29036 43372 29092 43374
rect 28924 43260 28980 43316
rect 29484 43820 29540 43876
rect 30044 44098 30100 44100
rect 30044 44046 30046 44098
rect 30046 44046 30098 44098
rect 30098 44046 30100 44098
rect 30044 44044 30100 44046
rect 29372 42812 29428 42868
rect 28588 42252 28644 42308
rect 28700 42028 28756 42084
rect 28028 40460 28084 40516
rect 28252 41356 28308 41412
rect 27916 40124 27972 40180
rect 27468 39340 27524 39396
rect 27804 38946 27860 38948
rect 27804 38894 27806 38946
rect 27806 38894 27858 38946
rect 27858 38894 27860 38946
rect 27804 38892 27860 38894
rect 27916 38780 27972 38836
rect 28028 39900 28084 39956
rect 27468 37772 27524 37828
rect 27804 37324 27860 37380
rect 27692 36764 27748 36820
rect 27468 35980 27524 36036
rect 28028 35980 28084 36036
rect 28140 39564 28196 39620
rect 27692 35868 27748 35924
rect 28588 41580 28644 41636
rect 28812 41468 28868 41524
rect 28924 42700 28980 42756
rect 28700 40012 28756 40068
rect 28476 39564 28532 39620
rect 28700 39394 28756 39396
rect 28700 39342 28702 39394
rect 28702 39342 28754 39394
rect 28754 39342 28756 39394
rect 28700 39340 28756 39342
rect 29148 41468 29204 41524
rect 29484 41916 29540 41972
rect 29260 40684 29316 40740
rect 29372 41244 29428 41300
rect 29372 40572 29428 40628
rect 30044 43596 30100 43652
rect 29820 43372 29876 43428
rect 29932 43260 29988 43316
rect 29708 42700 29764 42756
rect 29820 42812 29876 42868
rect 29820 42476 29876 42532
rect 30156 42866 30212 42868
rect 30156 42814 30158 42866
rect 30158 42814 30210 42866
rect 30210 42814 30212 42866
rect 30156 42812 30212 42814
rect 29932 42028 29988 42084
rect 29820 41970 29876 41972
rect 29820 41918 29822 41970
rect 29822 41918 29874 41970
rect 29874 41918 29876 41970
rect 29820 41916 29876 41918
rect 29596 41298 29652 41300
rect 29596 41246 29598 41298
rect 29598 41246 29650 41298
rect 29650 41246 29652 41298
rect 29596 41244 29652 41246
rect 29484 40684 29540 40740
rect 29708 40236 29764 40292
rect 30044 41468 30100 41524
rect 29820 40124 29876 40180
rect 29932 41020 29988 41076
rect 29820 39900 29876 39956
rect 28476 38834 28532 38836
rect 28476 38782 28478 38834
rect 28478 38782 28530 38834
rect 28530 38782 28532 38834
rect 28476 38780 28532 38782
rect 28700 38444 28756 38500
rect 28812 38892 28868 38948
rect 28924 37996 28980 38052
rect 28700 37826 28756 37828
rect 28700 37774 28702 37826
rect 28702 37774 28754 37826
rect 28754 37774 28756 37826
rect 28700 37772 28756 37774
rect 29372 39340 29428 39396
rect 29260 38946 29316 38948
rect 29260 38894 29262 38946
rect 29262 38894 29314 38946
rect 29314 38894 29316 38946
rect 29260 38892 29316 38894
rect 29820 39228 29876 39284
rect 30044 40460 30100 40516
rect 30828 47180 30884 47236
rect 31948 49196 32004 49252
rect 30940 45724 30996 45780
rect 31276 48636 31332 48692
rect 30828 45052 30884 45108
rect 31052 44994 31108 44996
rect 31052 44942 31054 44994
rect 31054 44942 31106 44994
rect 31106 44942 31108 44994
rect 31052 44940 31108 44942
rect 30940 44604 30996 44660
rect 31052 44716 31108 44772
rect 31836 48188 31892 48244
rect 31836 47404 31892 47460
rect 31948 47180 32004 47236
rect 31500 45778 31556 45780
rect 31500 45726 31502 45778
rect 31502 45726 31554 45778
rect 31554 45726 31556 45778
rect 31500 45724 31556 45726
rect 31500 45330 31556 45332
rect 31500 45278 31502 45330
rect 31502 45278 31554 45330
rect 31554 45278 31556 45330
rect 31500 45276 31556 45278
rect 32508 49756 32564 49812
rect 32396 48076 32452 48132
rect 32284 46508 32340 46564
rect 32172 45836 32228 45892
rect 32172 45612 32228 45668
rect 31164 44492 31220 44548
rect 31836 44492 31892 44548
rect 30380 43932 30436 43988
rect 30492 43708 30548 43764
rect 30380 42700 30436 42756
rect 30380 42476 30436 42532
rect 31724 44044 31780 44100
rect 30604 43596 30660 43652
rect 30380 41692 30436 41748
rect 30268 40908 30324 40964
rect 30380 41020 30436 41076
rect 30268 39788 30324 39844
rect 30716 41970 30772 41972
rect 30716 41918 30718 41970
rect 30718 41918 30770 41970
rect 30770 41918 30772 41970
rect 30716 41916 30772 41918
rect 30604 39676 30660 39732
rect 30940 43538 30996 43540
rect 30940 43486 30942 43538
rect 30942 43486 30994 43538
rect 30994 43486 30996 43538
rect 30940 43484 30996 43486
rect 31276 43538 31332 43540
rect 31276 43486 31278 43538
rect 31278 43486 31330 43538
rect 31330 43486 31332 43538
rect 31276 43484 31332 43486
rect 31500 43484 31556 43540
rect 31836 43484 31892 43540
rect 31276 42700 31332 42756
rect 31500 42700 31556 42756
rect 31388 42642 31444 42644
rect 31388 42590 31390 42642
rect 31390 42590 31442 42642
rect 31442 42590 31444 42642
rect 31388 42588 31444 42590
rect 31164 41804 31220 41860
rect 30828 41244 30884 41300
rect 30492 39394 30548 39396
rect 30492 39342 30494 39394
rect 30494 39342 30546 39394
rect 30546 39342 30548 39394
rect 30492 39340 30548 39342
rect 30940 40402 30996 40404
rect 30940 40350 30942 40402
rect 30942 40350 30994 40402
rect 30994 40350 30996 40402
rect 30940 40348 30996 40350
rect 31164 39730 31220 39732
rect 31164 39678 31166 39730
rect 31166 39678 31218 39730
rect 31218 39678 31220 39730
rect 31164 39676 31220 39678
rect 31612 42642 31668 42644
rect 31612 42590 31614 42642
rect 31614 42590 31666 42642
rect 31666 42590 31668 42642
rect 31612 42588 31668 42590
rect 31836 42588 31892 42644
rect 31388 41692 31444 41748
rect 32396 43708 32452 43764
rect 34972 49532 35028 49588
rect 34300 47292 34356 47348
rect 33068 47180 33124 47236
rect 33628 46060 33684 46116
rect 33628 45106 33684 45108
rect 33628 45054 33630 45106
rect 33630 45054 33682 45106
rect 33682 45054 33684 45106
rect 33628 45052 33684 45054
rect 32732 44098 32788 44100
rect 32732 44046 32734 44098
rect 32734 44046 32786 44098
rect 32786 44046 32788 44098
rect 32732 44044 32788 44046
rect 32508 43484 32564 43540
rect 31948 42252 32004 42308
rect 32396 43148 32452 43204
rect 31948 42082 32004 42084
rect 31948 42030 31950 42082
rect 31950 42030 32002 42082
rect 32002 42030 32004 42082
rect 31948 42028 32004 42030
rect 32172 42028 32228 42084
rect 31836 41916 31892 41972
rect 31500 40908 31556 40964
rect 31388 40460 31444 40516
rect 31388 40012 31444 40068
rect 31276 39116 31332 39172
rect 30492 38892 30548 38948
rect 31164 38892 31220 38948
rect 30380 38780 30436 38836
rect 30044 38556 30100 38612
rect 29708 38220 29764 38276
rect 29148 38108 29204 38164
rect 29484 38108 29540 38164
rect 28924 37826 28980 37828
rect 28924 37774 28926 37826
rect 28926 37774 28978 37826
rect 28978 37774 28980 37826
rect 28924 37772 28980 37774
rect 28588 37548 28644 37604
rect 29036 37548 29092 37604
rect 28364 36258 28420 36260
rect 28364 36206 28366 36258
rect 28366 36206 28418 36258
rect 28418 36206 28420 36258
rect 28364 36204 28420 36206
rect 28252 35980 28308 36036
rect 27132 35420 27188 35476
rect 26908 34300 26964 34356
rect 27020 34802 27076 34804
rect 27020 34750 27022 34802
rect 27022 34750 27074 34802
rect 27074 34750 27076 34802
rect 27020 34748 27076 34750
rect 26796 33964 26852 34020
rect 26908 33516 26964 33572
rect 26460 33122 26516 33124
rect 26460 33070 26462 33122
rect 26462 33070 26514 33122
rect 26514 33070 26516 33122
rect 26460 33068 26516 33070
rect 27132 34412 27188 34468
rect 27132 33628 27188 33684
rect 26124 31554 26180 31556
rect 26124 31502 26126 31554
rect 26126 31502 26178 31554
rect 26178 31502 26180 31554
rect 26124 31500 26180 31502
rect 26348 31500 26404 31556
rect 26124 31052 26180 31108
rect 26124 30882 26180 30884
rect 26124 30830 26126 30882
rect 26126 30830 26178 30882
rect 26178 30830 26180 30882
rect 26124 30828 26180 30830
rect 25116 30268 25172 30324
rect 24780 29986 24836 29988
rect 24780 29934 24782 29986
rect 24782 29934 24834 29986
rect 24834 29934 24836 29986
rect 24780 29932 24836 29934
rect 26572 32450 26628 32452
rect 26572 32398 26574 32450
rect 26574 32398 26626 32450
rect 26626 32398 26628 32450
rect 26572 32396 26628 32398
rect 27356 35532 27412 35588
rect 27692 35586 27748 35588
rect 27692 35534 27694 35586
rect 27694 35534 27746 35586
rect 27746 35534 27748 35586
rect 27692 35532 27748 35534
rect 27356 35084 27412 35140
rect 27580 35308 27636 35364
rect 27692 35196 27748 35252
rect 28588 36876 28644 36932
rect 28812 36204 28868 36260
rect 28588 35810 28644 35812
rect 28588 35758 28590 35810
rect 28590 35758 28642 35810
rect 28642 35758 28644 35810
rect 28588 35756 28644 35758
rect 29484 37772 29540 37828
rect 29260 37378 29316 37380
rect 29260 37326 29262 37378
rect 29262 37326 29314 37378
rect 29314 37326 29316 37378
rect 29260 37324 29316 37326
rect 28476 35196 28532 35252
rect 29260 36204 29316 36260
rect 27580 34412 27636 34468
rect 27468 33458 27524 33460
rect 27468 33406 27470 33458
rect 27470 33406 27522 33458
rect 27522 33406 27524 33458
rect 27468 33404 27524 33406
rect 27468 32956 27524 33012
rect 27244 32508 27300 32564
rect 26572 31778 26628 31780
rect 26572 31726 26574 31778
rect 26574 31726 26626 31778
rect 26626 31726 26628 31778
rect 26572 31724 26628 31726
rect 26572 31388 26628 31444
rect 26796 31500 26852 31556
rect 26796 31164 26852 31220
rect 27916 34636 27972 34692
rect 28028 34354 28084 34356
rect 28028 34302 28030 34354
rect 28030 34302 28082 34354
rect 28082 34302 28084 34354
rect 28028 34300 28084 34302
rect 28028 33852 28084 33908
rect 28588 34914 28644 34916
rect 28588 34862 28590 34914
rect 28590 34862 28642 34914
rect 28642 34862 28644 34914
rect 28588 34860 28644 34862
rect 28140 33404 28196 33460
rect 28476 34412 28532 34468
rect 29148 35922 29204 35924
rect 29148 35870 29150 35922
rect 29150 35870 29202 35922
rect 29202 35870 29204 35922
rect 29148 35868 29204 35870
rect 29596 37938 29652 37940
rect 29596 37886 29598 37938
rect 29598 37886 29650 37938
rect 29650 37886 29652 37938
rect 29596 37884 29652 37886
rect 29708 37772 29764 37828
rect 29708 37548 29764 37604
rect 29596 37436 29652 37492
rect 29708 37266 29764 37268
rect 29708 37214 29710 37266
rect 29710 37214 29762 37266
rect 29762 37214 29764 37266
rect 29708 37212 29764 37214
rect 30268 38332 30324 38388
rect 30156 38274 30212 38276
rect 30156 38222 30158 38274
rect 30158 38222 30210 38274
rect 30210 38222 30212 38274
rect 30156 38220 30212 38222
rect 31052 38444 31108 38500
rect 30044 37772 30100 37828
rect 30044 37212 30100 37268
rect 29820 36988 29876 37044
rect 29932 36540 29988 36596
rect 30156 36540 30212 36596
rect 29036 33852 29092 33908
rect 29596 35756 29652 35812
rect 30380 37378 30436 37380
rect 30380 37326 30382 37378
rect 30382 37326 30434 37378
rect 30434 37326 30436 37378
rect 30380 37324 30436 37326
rect 30380 36706 30436 36708
rect 30380 36654 30382 36706
rect 30382 36654 30434 36706
rect 30434 36654 30436 36706
rect 30380 36652 30436 36654
rect 30828 37826 30884 37828
rect 30828 37774 30830 37826
rect 30830 37774 30882 37826
rect 30882 37774 30884 37826
rect 30828 37772 30884 37774
rect 30716 36652 30772 36708
rect 30380 36482 30436 36484
rect 30380 36430 30382 36482
rect 30382 36430 30434 36482
rect 30434 36430 30436 36482
rect 30380 36428 30436 36430
rect 30604 36092 30660 36148
rect 28924 33628 28980 33684
rect 28812 33458 28868 33460
rect 28812 33406 28814 33458
rect 28814 33406 28866 33458
rect 28866 33406 28868 33458
rect 28812 33404 28868 33406
rect 28700 33180 28756 33236
rect 28476 33068 28532 33124
rect 28364 32844 28420 32900
rect 29484 35308 29540 35364
rect 29708 35420 29764 35476
rect 29820 35532 29876 35588
rect 29372 34130 29428 34132
rect 29372 34078 29374 34130
rect 29374 34078 29426 34130
rect 29426 34078 29428 34130
rect 29372 34076 29428 34078
rect 29484 33628 29540 33684
rect 29260 32956 29316 33012
rect 28476 32284 28532 32340
rect 30156 35308 30212 35364
rect 29932 35084 29988 35140
rect 30940 37100 30996 37156
rect 30828 36540 30884 36596
rect 30492 34914 30548 34916
rect 30492 34862 30494 34914
rect 30494 34862 30546 34914
rect 30546 34862 30548 34914
rect 30492 34860 30548 34862
rect 29820 34188 29876 34244
rect 29708 32172 29764 32228
rect 28252 30380 28308 30436
rect 27804 29820 27860 29876
rect 26460 27916 26516 27972
rect 28588 28140 28644 28196
rect 28588 26348 28644 26404
rect 30380 34524 30436 34580
rect 30156 34188 30212 34244
rect 30044 27468 30100 27524
rect 30268 31612 30324 31668
rect 29932 26236 29988 26292
rect 30828 35308 30884 35364
rect 30940 35196 30996 35252
rect 30940 35026 30996 35028
rect 30940 34974 30942 35026
rect 30942 34974 30994 35026
rect 30994 34974 30996 35026
rect 30940 34972 30996 34974
rect 30716 34354 30772 34356
rect 30716 34302 30718 34354
rect 30718 34302 30770 34354
rect 30770 34302 30772 34354
rect 30716 34300 30772 34302
rect 31276 38444 31332 38500
rect 31276 38220 31332 38276
rect 31276 37772 31332 37828
rect 31500 37996 31556 38052
rect 31500 37436 31556 37492
rect 32060 41580 32116 41636
rect 32284 40908 32340 40964
rect 33068 43372 33124 43428
rect 32732 42924 32788 42980
rect 32508 42530 32564 42532
rect 32508 42478 32510 42530
rect 32510 42478 32562 42530
rect 32562 42478 32564 42530
rect 32508 42476 32564 42478
rect 33068 42642 33124 42644
rect 33068 42590 33070 42642
rect 33070 42590 33122 42642
rect 33122 42590 33124 42642
rect 33068 42588 33124 42590
rect 32844 42140 32900 42196
rect 32620 41804 32676 41860
rect 32508 41580 32564 41636
rect 32396 41186 32452 41188
rect 32396 41134 32398 41186
rect 32398 41134 32450 41186
rect 32450 41134 32452 41186
rect 32396 41132 32452 41134
rect 32284 40460 32340 40516
rect 32060 40178 32116 40180
rect 32060 40126 32062 40178
rect 32062 40126 32114 40178
rect 32114 40126 32116 40178
rect 32060 40124 32116 40126
rect 31948 39676 32004 39732
rect 31724 39340 31780 39396
rect 33516 43148 33572 43204
rect 33516 42924 33572 42980
rect 33180 41356 33236 41412
rect 33292 42588 33348 42644
rect 33852 45948 33908 46004
rect 33740 44604 33796 44660
rect 33740 43148 33796 43204
rect 34076 43036 34132 43092
rect 33292 41692 33348 41748
rect 33068 41186 33124 41188
rect 33068 41134 33070 41186
rect 33070 41134 33122 41186
rect 33122 41134 33124 41186
rect 33068 41132 33124 41134
rect 33404 41580 33460 41636
rect 33516 41692 33572 41748
rect 33404 41132 33460 41188
rect 32620 40908 32676 40964
rect 33180 40962 33236 40964
rect 33180 40910 33182 40962
rect 33182 40910 33234 40962
rect 33234 40910 33236 40962
rect 33180 40908 33236 40910
rect 33964 42476 34020 42532
rect 34860 45218 34916 45220
rect 34860 45166 34862 45218
rect 34862 45166 34914 45218
rect 34914 45166 34916 45218
rect 34860 45164 34916 45166
rect 34524 44098 34580 44100
rect 34524 44046 34526 44098
rect 34526 44046 34578 44098
rect 34578 44046 34580 44098
rect 34524 44044 34580 44046
rect 34412 43820 34468 43876
rect 34972 43932 35028 43988
rect 34860 43820 34916 43876
rect 34748 43484 34804 43540
rect 34748 43148 34804 43204
rect 34860 43036 34916 43092
rect 34524 42978 34580 42980
rect 34524 42926 34526 42978
rect 34526 42926 34578 42978
rect 34578 42926 34580 42978
rect 34524 42924 34580 42926
rect 34972 42588 35028 42644
rect 33852 41020 33908 41076
rect 33628 40908 33684 40964
rect 33404 40572 33460 40628
rect 33628 40572 33684 40628
rect 32732 40460 32788 40516
rect 32956 40460 33012 40516
rect 32620 40402 32676 40404
rect 32620 40350 32622 40402
rect 32622 40350 32674 40402
rect 32674 40350 32676 40402
rect 32620 40348 32676 40350
rect 33964 40402 34020 40404
rect 33964 40350 33966 40402
rect 33966 40350 34018 40402
rect 34018 40350 34020 40402
rect 33964 40348 34020 40350
rect 32508 40178 32564 40180
rect 32508 40126 32510 40178
rect 32510 40126 32562 40178
rect 32562 40126 32564 40178
rect 32508 40124 32564 40126
rect 32508 39900 32564 39956
rect 33068 40012 33124 40068
rect 32396 39116 32452 39172
rect 32732 39676 32788 39732
rect 32172 38946 32228 38948
rect 32172 38894 32174 38946
rect 32174 38894 32226 38946
rect 32226 38894 32228 38946
rect 32172 38892 32228 38894
rect 32396 38834 32452 38836
rect 32396 38782 32398 38834
rect 32398 38782 32450 38834
rect 32450 38782 32452 38834
rect 32396 38780 32452 38782
rect 31948 38722 32004 38724
rect 31948 38670 31950 38722
rect 31950 38670 32002 38722
rect 32002 38670 32004 38722
rect 31948 38668 32004 38670
rect 33180 39676 33236 39732
rect 31724 38444 31780 38500
rect 31948 38444 32004 38500
rect 31836 38332 31892 38388
rect 31724 36876 31780 36932
rect 31612 36652 31668 36708
rect 31724 36370 31780 36372
rect 31724 36318 31726 36370
rect 31726 36318 31778 36370
rect 31778 36318 31780 36370
rect 31724 36316 31780 36318
rect 31276 36092 31332 36148
rect 31276 35868 31332 35924
rect 31164 35196 31220 35252
rect 31164 33628 31220 33684
rect 31612 36204 31668 36260
rect 31612 35868 31668 35924
rect 31500 35698 31556 35700
rect 31500 35646 31502 35698
rect 31502 35646 31554 35698
rect 31554 35646 31556 35698
rect 31500 35644 31556 35646
rect 32844 39116 32900 39172
rect 32732 39004 32788 39060
rect 31948 36316 32004 36372
rect 31948 35922 32004 35924
rect 31948 35870 31950 35922
rect 31950 35870 32002 35922
rect 32002 35870 32004 35922
rect 31948 35868 32004 35870
rect 31276 33852 31332 33908
rect 31276 33516 31332 33572
rect 31052 32732 31108 32788
rect 31948 33404 32004 33460
rect 30604 29484 30660 29540
rect 30268 24668 30324 24724
rect 32172 37154 32228 37156
rect 32172 37102 32174 37154
rect 32174 37102 32226 37154
rect 32226 37102 32228 37154
rect 32172 37100 32228 37102
rect 32172 36540 32228 36596
rect 32172 36092 32228 36148
rect 32396 35810 32452 35812
rect 32396 35758 32398 35810
rect 32398 35758 32450 35810
rect 32450 35758 32452 35810
rect 32396 35756 32452 35758
rect 32284 34860 32340 34916
rect 32172 34690 32228 34692
rect 32172 34638 32174 34690
rect 32174 34638 32226 34690
rect 32226 34638 32228 34690
rect 32172 34636 32228 34638
rect 32172 34076 32228 34132
rect 32620 38050 32676 38052
rect 32620 37998 32622 38050
rect 32622 37998 32674 38050
rect 32674 37998 32676 38050
rect 32620 37996 32676 37998
rect 33068 38780 33124 38836
rect 33292 39228 33348 39284
rect 33628 39618 33684 39620
rect 33628 39566 33630 39618
rect 33630 39566 33682 39618
rect 33682 39566 33684 39618
rect 33628 39564 33684 39566
rect 33516 39228 33572 39284
rect 33740 39228 33796 39284
rect 33852 39564 33908 39620
rect 33404 39004 33460 39060
rect 33516 38780 33572 38836
rect 33964 38834 34020 38836
rect 33964 38782 33966 38834
rect 33966 38782 34018 38834
rect 34018 38782 34020 38834
rect 33964 38780 34020 38782
rect 33516 37660 33572 37716
rect 34972 42364 35028 42420
rect 34636 41580 34692 41636
rect 34748 42028 34804 42084
rect 34188 41468 34244 41524
rect 34636 41356 34692 41412
rect 34412 41298 34468 41300
rect 34412 41246 34414 41298
rect 34414 41246 34466 41298
rect 34466 41246 34468 41298
rect 34412 41244 34468 41246
rect 34300 40684 34356 40740
rect 34188 40402 34244 40404
rect 34188 40350 34190 40402
rect 34190 40350 34242 40402
rect 34242 40350 34244 40402
rect 34188 40348 34244 40350
rect 38332 49308 38388 49364
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 37324 48972 37380 49028
rect 36988 48748 37044 48804
rect 35868 47740 35924 47796
rect 35644 45500 35700 45556
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35308 44492 35364 44548
rect 35532 44380 35588 44436
rect 35308 44210 35364 44212
rect 35308 44158 35310 44210
rect 35310 44158 35362 44210
rect 35362 44158 35364 44210
rect 35308 44156 35364 44158
rect 35756 44380 35812 44436
rect 35756 43596 35812 43652
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35756 43148 35812 43204
rect 35532 42924 35588 42980
rect 35252 42812 35308 42868
rect 35644 42700 35700 42756
rect 36316 47516 36372 47572
rect 36204 47068 36260 47124
rect 36092 45890 36148 45892
rect 36092 45838 36094 45890
rect 36094 45838 36146 45890
rect 36146 45838 36148 45890
rect 36092 45836 36148 45838
rect 35308 41916 35364 41972
rect 35084 41746 35140 41748
rect 35084 41694 35086 41746
rect 35086 41694 35138 41746
rect 35138 41694 35140 41746
rect 35084 41692 35140 41694
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35644 41468 35700 41524
rect 34972 41132 35028 41188
rect 35196 41244 35252 41300
rect 34860 40684 34916 40740
rect 34636 40012 34692 40068
rect 34300 39228 34356 39284
rect 34412 39900 34468 39956
rect 34972 40908 35028 40964
rect 34076 38556 34132 38612
rect 34188 38892 34244 38948
rect 34524 38332 34580 38388
rect 33964 37938 34020 37940
rect 33964 37886 33966 37938
rect 33966 37886 34018 37938
rect 34018 37886 34020 37938
rect 33964 37884 34020 37886
rect 33740 37660 33796 37716
rect 33964 37378 34020 37380
rect 33964 37326 33966 37378
rect 33966 37326 34018 37378
rect 34018 37326 34020 37378
rect 33964 37324 34020 37326
rect 33516 37266 33572 37268
rect 33516 37214 33518 37266
rect 33518 37214 33570 37266
rect 33570 37214 33572 37266
rect 33516 37212 33572 37214
rect 32956 36988 33012 37044
rect 32508 31276 32564 31332
rect 32620 36876 32676 36932
rect 32732 36764 32788 36820
rect 32844 36204 32900 36260
rect 32732 36092 32788 36148
rect 32732 35196 32788 35252
rect 32732 33404 32788 33460
rect 32844 31724 32900 31780
rect 32620 28700 32676 28756
rect 34636 37996 34692 38052
rect 33516 36316 33572 36372
rect 33068 35980 33124 36036
rect 34524 37324 34580 37380
rect 34412 37154 34468 37156
rect 34412 37102 34414 37154
rect 34414 37102 34466 37154
rect 34466 37102 34468 37154
rect 34412 37100 34468 37102
rect 33628 35644 33684 35700
rect 32956 28028 33012 28084
rect 33852 33292 33908 33348
rect 34412 32956 34468 33012
rect 34748 39340 34804 39396
rect 34748 39116 34804 39172
rect 36204 43036 36260 43092
rect 37100 45666 37156 45668
rect 37100 45614 37102 45666
rect 37102 45614 37154 45666
rect 37154 45614 37156 45666
rect 37100 45612 37156 45614
rect 37212 45388 37268 45444
rect 36652 44098 36708 44100
rect 36652 44046 36654 44098
rect 36654 44046 36706 44098
rect 36706 44046 36708 44098
rect 36652 44044 36708 44046
rect 36652 43260 36708 43316
rect 36652 42754 36708 42756
rect 36652 42702 36654 42754
rect 36654 42702 36706 42754
rect 36706 42702 36708 42754
rect 36652 42700 36708 42702
rect 36876 43820 36932 43876
rect 36876 43148 36932 43204
rect 36764 41916 36820 41972
rect 35532 40962 35588 40964
rect 35532 40910 35534 40962
rect 35534 40910 35586 40962
rect 35586 40910 35588 40962
rect 35532 40908 35588 40910
rect 35196 40684 35252 40740
rect 35420 40796 35476 40852
rect 35644 40796 35700 40852
rect 35644 40348 35700 40404
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35084 39788 35140 39844
rect 35084 39506 35140 39508
rect 35084 39454 35086 39506
rect 35086 39454 35138 39506
rect 35138 39454 35140 39506
rect 35084 39452 35140 39454
rect 35308 39788 35364 39844
rect 35756 39900 35812 39956
rect 35196 39228 35252 39284
rect 35420 39116 35476 39172
rect 35532 39004 35588 39060
rect 35084 38780 35140 38836
rect 35308 38834 35364 38836
rect 35308 38782 35310 38834
rect 35310 38782 35362 38834
rect 35362 38782 35364 38834
rect 35308 38780 35364 38782
rect 36092 41244 36148 41300
rect 36428 40962 36484 40964
rect 36428 40910 36430 40962
rect 36430 40910 36482 40962
rect 36482 40910 36484 40962
rect 36428 40908 36484 40910
rect 36428 40402 36484 40404
rect 36428 40350 36430 40402
rect 36430 40350 36482 40402
rect 36482 40350 36484 40402
rect 36428 40348 36484 40350
rect 34860 38108 34916 38164
rect 34860 37884 34916 37940
rect 34860 37490 34916 37492
rect 34860 37438 34862 37490
rect 34862 37438 34914 37490
rect 34914 37438 34916 37490
rect 34860 37436 34916 37438
rect 34972 34636 35028 34692
rect 34748 31164 34804 31220
rect 34524 29708 34580 29764
rect 36092 39340 36148 39396
rect 36204 39058 36260 39060
rect 36204 39006 36206 39058
rect 36206 39006 36258 39058
rect 36258 39006 36260 39058
rect 36204 39004 36260 39006
rect 36316 38892 36372 38948
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35980 38556 36036 38612
rect 36092 38668 36148 38724
rect 35868 38444 35924 38500
rect 35756 38050 35812 38052
rect 35756 37998 35758 38050
rect 35758 37998 35810 38050
rect 35810 37998 35812 38050
rect 35756 37996 35812 37998
rect 35308 37826 35364 37828
rect 35308 37774 35310 37826
rect 35310 37774 35362 37826
rect 35362 37774 35364 37826
rect 35308 37772 35364 37774
rect 35756 37772 35812 37828
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35644 36092 35700 36148
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35868 34524 35924 34580
rect 35532 34412 35588 34468
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 36428 37548 36484 37604
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35084 29260 35140 29316
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 33852 26796 33908 26852
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 32060 23996 32116 24052
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 31948 18284 32004 18340
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 36092 32508 36148 32564
rect 36652 41186 36708 41188
rect 36652 41134 36654 41186
rect 36654 41134 36706 41186
rect 36706 41134 36708 41186
rect 36652 41132 36708 41134
rect 36652 39116 36708 39172
rect 36652 30940 36708 30996
rect 36876 37212 36932 37268
rect 37436 47628 37492 47684
rect 37548 46396 37604 46452
rect 38444 49084 38500 49140
rect 39228 48524 39284 48580
rect 38892 47852 38948 47908
rect 39452 48188 39508 48244
rect 39340 46396 39396 46452
rect 37548 44994 37604 44996
rect 37548 44942 37550 44994
rect 37550 44942 37602 44994
rect 37602 44942 37604 44994
rect 37548 44940 37604 44942
rect 37548 43260 37604 43316
rect 37436 41804 37492 41860
rect 37436 40962 37492 40964
rect 37436 40910 37438 40962
rect 37438 40910 37490 40962
rect 37490 40910 37492 40962
rect 37436 40908 37492 40910
rect 38220 45052 38276 45108
rect 37772 44828 37828 44884
rect 37884 43820 37940 43876
rect 38108 43708 38164 43764
rect 37996 43538 38052 43540
rect 37996 43486 37998 43538
rect 37998 43486 38050 43538
rect 38050 43486 38052 43538
rect 37996 43484 38052 43486
rect 38108 42476 38164 42532
rect 38332 44828 38388 44884
rect 38780 44322 38836 44324
rect 38780 44270 38782 44322
rect 38782 44270 38834 44322
rect 38834 44270 38836 44322
rect 38780 44268 38836 44270
rect 38332 44156 38388 44212
rect 38332 43708 38388 43764
rect 38668 44156 38724 44212
rect 38892 43762 38948 43764
rect 38892 43710 38894 43762
rect 38894 43710 38946 43762
rect 38946 43710 38948 43762
rect 38892 43708 38948 43710
rect 39564 47516 39620 47572
rect 40684 48300 40740 48356
rect 40348 47068 40404 47124
rect 38444 42028 38500 42084
rect 38332 41074 38388 41076
rect 38332 41022 38334 41074
rect 38334 41022 38386 41074
rect 38386 41022 38388 41074
rect 38332 41020 38388 41022
rect 37884 40962 37940 40964
rect 37884 40910 37886 40962
rect 37886 40910 37938 40962
rect 37938 40910 37940 40962
rect 37884 40908 37940 40910
rect 37884 40684 37940 40740
rect 38220 40626 38276 40628
rect 38220 40574 38222 40626
rect 38222 40574 38274 40626
rect 38274 40574 38276 40626
rect 38220 40572 38276 40574
rect 37100 39900 37156 39956
rect 37548 38946 37604 38948
rect 37548 38894 37550 38946
rect 37550 38894 37602 38946
rect 37602 38894 37604 38946
rect 37548 38892 37604 38894
rect 37324 38444 37380 38500
rect 36988 33068 37044 33124
rect 37884 40236 37940 40292
rect 38332 39618 38388 39620
rect 38332 39566 38334 39618
rect 38334 39566 38386 39618
rect 38386 39566 38388 39618
rect 38332 39564 38388 39566
rect 38668 42476 38724 42532
rect 38668 40460 38724 40516
rect 38668 40290 38724 40292
rect 38668 40238 38670 40290
rect 38670 40238 38722 40290
rect 38722 40238 38724 40290
rect 38668 40236 38724 40238
rect 38780 39618 38836 39620
rect 38780 39566 38782 39618
rect 38782 39566 38834 39618
rect 38834 39566 38836 39618
rect 38780 39564 38836 39566
rect 39228 43596 39284 43652
rect 39676 43484 39732 43540
rect 39900 43820 39956 43876
rect 39788 43426 39844 43428
rect 39788 43374 39790 43426
rect 39790 43374 39842 43426
rect 39842 43374 39844 43426
rect 39788 43372 39844 43374
rect 39228 42530 39284 42532
rect 39228 42478 39230 42530
rect 39230 42478 39282 42530
rect 39282 42478 39284 42530
rect 39228 42476 39284 42478
rect 39340 42812 39396 42868
rect 39116 41858 39172 41860
rect 39116 41806 39118 41858
rect 39118 41806 39170 41858
rect 39170 41806 39172 41858
rect 39116 41804 39172 41806
rect 39228 40962 39284 40964
rect 39228 40910 39230 40962
rect 39230 40910 39282 40962
rect 39282 40910 39284 40962
rect 39228 40908 39284 40910
rect 39116 40402 39172 40404
rect 39116 40350 39118 40402
rect 39118 40350 39170 40402
rect 39170 40350 39172 40402
rect 39116 40348 39172 40350
rect 39452 38556 39508 38612
rect 39564 37996 39620 38052
rect 39340 36540 39396 36596
rect 39004 35532 39060 35588
rect 38556 35084 38612 35140
rect 37996 32508 38052 32564
rect 40124 42812 40180 42868
rect 40124 42642 40180 42644
rect 40124 42590 40126 42642
rect 40126 42590 40178 42642
rect 40178 42590 40180 42642
rect 40124 42588 40180 42590
rect 40124 41074 40180 41076
rect 40124 41022 40126 41074
rect 40126 41022 40178 41074
rect 40178 41022 40180 41074
rect 40124 41020 40180 41022
rect 40012 38780 40068 38836
rect 40236 33964 40292 34020
rect 37660 31836 37716 31892
rect 36764 30828 36820 30884
rect 36540 29596 36596 29652
rect 36092 16716 36148 16772
rect 37212 26796 37268 26852
rect 35644 15036 35700 15092
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 23772 11676 23828 11732
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 19628 11340 19684 11396
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 36428 3442 36484 3444
rect 36428 3390 36430 3442
rect 36430 3390 36482 3442
rect 36482 3390 36484 3442
rect 36428 3388 36484 3390
rect 36988 3388 37044 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 28252 3276 28308 3332
rect 29260 3330 29316 3332
rect 29260 3278 29262 3330
rect 29262 3278 29314 3330
rect 29314 3278 29316 3330
rect 29260 3276 29316 3278
rect 40572 45612 40628 45668
rect 41804 45890 41860 45892
rect 41804 45838 41806 45890
rect 41806 45838 41858 45890
rect 41858 45838 41860 45890
rect 41804 45836 41860 45838
rect 41356 45778 41412 45780
rect 41356 45726 41358 45778
rect 41358 45726 41410 45778
rect 41410 45726 41412 45778
rect 41356 45724 41412 45726
rect 40908 45666 40964 45668
rect 40908 45614 40910 45666
rect 40910 45614 40962 45666
rect 40962 45614 40964 45666
rect 40908 45612 40964 45614
rect 40572 42364 40628 42420
rect 40460 41692 40516 41748
rect 40572 41356 40628 41412
rect 47740 45612 47796 45668
rect 47292 43036 47348 43092
rect 48076 43036 48132 43092
rect 41468 40012 41524 40068
rect 42028 41580 42084 41636
rect 40908 39004 40964 39060
rect 40348 21756 40404 21812
rect 40012 19852 40068 19908
rect 48076 39676 48132 39732
rect 48076 37660 48132 37716
rect 48076 35644 48132 35700
rect 48076 34300 48132 34356
rect 42028 18396 42084 18452
rect 47740 33852 47796 33908
rect 37548 3442 37604 3444
rect 37548 3390 37550 3442
rect 37550 3390 37602 3442
rect 37602 3390 37604 3442
rect 37548 3388 37604 3390
rect 47516 3388 47572 3444
rect 48076 32284 48132 32340
rect 48076 30940 48132 30996
rect 48076 28924 48132 28980
rect 48076 26850 48132 26852
rect 48076 26798 48078 26850
rect 48078 26798 48130 26850
rect 48130 26798 48132 26850
rect 48076 26796 48132 26798
rect 48076 23548 48132 23604
rect 48076 21532 48132 21588
rect 48076 18562 48132 18564
rect 48076 18510 48078 18562
rect 48078 18510 48130 18562
rect 48130 18510 48132 18562
rect 48076 18508 48132 18510
rect 48076 16828 48132 16884
rect 48076 12850 48132 12852
rect 48076 12798 48078 12850
rect 48078 12798 48130 12850
rect 48130 12798 48132 12850
rect 48076 12796 48132 12798
rect 48076 11452 48132 11508
rect 48076 9436 48132 9492
rect 48076 7420 48132 7476
rect 48076 6076 48132 6132
rect 48076 3442 48132 3444
rect 48076 3390 48078 3442
rect 48078 3390 48130 3442
rect 48130 3390 48132 3442
rect 48076 3388 48132 3390
rect 48188 2044 48244 2100
rect 49084 3388 49140 3444
rect 47180 700 47236 756
<< metal3 >>
rect 3266 49868 3276 49924
rect 3332 49868 12236 49924
rect 12292 49868 12302 49924
rect 21522 49868 21532 49924
rect 21588 49868 32060 49924
rect 32116 49868 32126 49924
rect 32284 49868 34748 49924
rect 34804 49868 34814 49924
rect 32284 49812 32340 49868
rect 11666 49756 11676 49812
rect 11732 49756 25788 49812
rect 25844 49756 25854 49812
rect 26114 49756 26124 49812
rect 26180 49756 32340 49812
rect 32498 49756 32508 49812
rect 32564 49756 32574 49812
rect 32508 49700 32564 49756
rect 10658 49644 10668 49700
rect 10724 49644 24892 49700
rect 24948 49644 24958 49700
rect 25778 49644 25788 49700
rect 25844 49644 32564 49700
rect 8082 49532 8092 49588
rect 8148 49532 17948 49588
rect 18004 49532 18014 49588
rect 18946 49532 18956 49588
rect 19012 49532 26012 49588
rect 26068 49532 26078 49588
rect 26226 49532 26236 49588
rect 26292 49532 34972 49588
rect 35028 49532 35038 49588
rect 9538 49420 9548 49476
rect 9604 49420 25788 49476
rect 25844 49420 25854 49476
rect 26002 49420 26012 49476
rect 26068 49420 30492 49476
rect 30548 49420 30558 49476
rect 6972 49308 16828 49364
rect 16884 49308 16894 49364
rect 23202 49308 23212 49364
rect 23268 49308 26348 49364
rect 26404 49308 26414 49364
rect 26572 49308 38332 49364
rect 38388 49308 38398 49364
rect 6972 49252 7028 49308
rect 26572 49252 26628 49308
rect 6962 49196 6972 49252
rect 7028 49196 7038 49252
rect 11666 49196 11676 49252
rect 11732 49196 26012 49252
rect 26068 49196 26078 49252
rect 26562 49196 26572 49252
rect 26628 49196 26638 49252
rect 26786 49196 26796 49252
rect 26852 49196 31948 49252
rect 32004 49196 32014 49252
rect 200 49140 800 49168
rect 200 49084 3164 49140
rect 3220 49084 3230 49140
rect 11554 49084 11564 49140
rect 11620 49084 15708 49140
rect 15764 49084 15774 49140
rect 18050 49084 18060 49140
rect 18116 49084 26012 49140
rect 26068 49084 26078 49140
rect 26236 49084 38444 49140
rect 38500 49084 38510 49140
rect 200 49056 800 49084
rect 26236 49028 26292 49084
rect 5170 48972 5180 49028
rect 5236 48972 13804 49028
rect 13860 48972 13870 49028
rect 16818 48972 16828 49028
rect 16884 48972 18284 49028
rect 18340 48972 18350 49028
rect 22754 48972 22764 49028
rect 22820 48972 25564 49028
rect 25620 48972 25630 49028
rect 25778 48972 25788 49028
rect 25844 48972 26292 49028
rect 26450 48972 26460 49028
rect 26516 48972 37324 49028
rect 37380 48972 37390 49028
rect 5954 48860 5964 48916
rect 6020 48860 8428 48916
rect 10770 48860 10780 48916
rect 10836 48860 27804 48916
rect 27860 48860 27870 48916
rect 8372 48804 8428 48860
rect 8372 48748 14588 48804
rect 14644 48748 14654 48804
rect 14802 48748 14812 48804
rect 14868 48748 22988 48804
rect 23044 48748 23054 48804
rect 26002 48748 26012 48804
rect 26068 48748 36988 48804
rect 37044 48748 37054 48804
rect 4946 48636 4956 48692
rect 5012 48636 16492 48692
rect 16548 48636 16558 48692
rect 18946 48636 18956 48692
rect 19012 48636 25788 48692
rect 25844 48636 25854 48692
rect 26460 48636 26908 48692
rect 27010 48636 27020 48692
rect 27076 48636 31276 48692
rect 31332 48636 31342 48692
rect 26460 48580 26516 48636
rect 8372 48524 16604 48580
rect 16660 48524 16670 48580
rect 16930 48524 16940 48580
rect 16996 48524 26516 48580
rect 26852 48580 26908 48636
rect 26852 48524 29036 48580
rect 29092 48524 29102 48580
rect 30146 48524 30156 48580
rect 30212 48524 39228 48580
rect 39284 48524 39294 48580
rect 8372 48356 8428 48524
rect 11106 48412 11116 48468
rect 11172 48412 14812 48468
rect 14868 48412 14878 48468
rect 16930 48412 16940 48468
rect 16996 48412 26796 48468
rect 26852 48412 26862 48468
rect 27346 48412 27356 48468
rect 27412 48412 30604 48468
rect 30660 48412 30670 48468
rect 30818 48412 30828 48468
rect 30884 48412 38668 48468
rect 38612 48356 38668 48412
rect 49200 48384 49800 48496
rect 2258 48300 2268 48356
rect 2324 48300 8428 48356
rect 9314 48300 9324 48356
rect 9380 48300 28812 48356
rect 28868 48300 28878 48356
rect 29362 48300 29372 48356
rect 29428 48300 36316 48356
rect 36372 48300 36382 48356
rect 38612 48300 40684 48356
rect 40740 48300 40750 48356
rect 7970 48188 7980 48244
rect 8036 48188 30380 48244
rect 30436 48188 30446 48244
rect 31826 48188 31836 48244
rect 31892 48188 39452 48244
rect 39508 48188 39518 48244
rect 5058 48076 5068 48132
rect 5124 48076 11620 48132
rect 11778 48076 11788 48132
rect 11844 48076 32396 48132
rect 32452 48076 32462 48132
rect 11564 48020 11620 48076
rect 3826 47964 3836 48020
rect 3892 47964 8372 48020
rect 8428 47964 8438 48020
rect 8530 47964 8540 48020
rect 8596 47964 11340 48020
rect 11396 47964 11406 48020
rect 11564 47964 13468 48020
rect 13524 47964 13534 48020
rect 14018 47964 14028 48020
rect 14084 47964 26572 48020
rect 26628 47964 26638 48020
rect 27010 47964 27020 48020
rect 27076 47964 34300 48020
rect 34356 47964 34366 48020
rect 7858 47852 7868 47908
rect 7924 47852 15596 47908
rect 15652 47852 15662 47908
rect 15810 47852 15820 47908
rect 15876 47852 29596 47908
rect 29652 47852 29662 47908
rect 29810 47852 29820 47908
rect 29876 47852 38892 47908
rect 38948 47852 38958 47908
rect 200 47796 800 47824
rect 200 47740 1820 47796
rect 1876 47740 1886 47796
rect 6850 47740 6860 47796
rect 6916 47740 8428 47796
rect 8484 47740 8494 47796
rect 8754 47740 8764 47796
rect 8820 47740 16940 47796
rect 16996 47740 17006 47796
rect 17826 47740 17836 47796
rect 17892 47740 28924 47796
rect 28980 47740 30156 47796
rect 30212 47740 30222 47796
rect 30594 47740 30604 47796
rect 30660 47740 35868 47796
rect 35924 47740 35934 47796
rect 200 47712 800 47740
rect 6066 47628 6076 47684
rect 6132 47628 8316 47684
rect 8372 47628 8596 47684
rect 10546 47628 10556 47684
rect 10612 47628 14700 47684
rect 14756 47628 14766 47684
rect 14914 47628 14924 47684
rect 14980 47628 27804 47684
rect 27860 47628 27870 47684
rect 29474 47628 29484 47684
rect 29540 47628 37436 47684
rect 37492 47628 37502 47684
rect 8540 47572 8596 47628
rect 7074 47516 7084 47572
rect 7140 47516 8428 47572
rect 8540 47516 16716 47572
rect 16772 47516 16782 47572
rect 16930 47516 16940 47572
rect 16996 47516 25452 47572
rect 25508 47516 25518 47572
rect 27234 47516 27244 47572
rect 27300 47516 36316 47572
rect 36372 47516 36382 47572
rect 38612 47516 39564 47572
rect 39620 47516 39630 47572
rect 8372 47460 8428 47516
rect 38612 47460 38668 47516
rect 8372 47404 13916 47460
rect 13972 47404 13982 47460
rect 14130 47404 14140 47460
rect 14196 47404 23156 47460
rect 23314 47404 23324 47460
rect 23380 47404 30716 47460
rect 30772 47404 31836 47460
rect 31892 47404 31902 47460
rect 36306 47404 36316 47460
rect 36372 47404 38668 47460
rect 23100 47348 23156 47404
rect 690 47292 700 47348
rect 756 47292 2492 47348
rect 2548 47292 2558 47348
rect 9090 47292 9100 47348
rect 9156 47292 18508 47348
rect 18564 47292 20188 47348
rect 23100 47292 23660 47348
rect 23716 47292 23726 47348
rect 23874 47292 23884 47348
rect 23940 47292 27356 47348
rect 27412 47292 27422 47348
rect 27570 47292 27580 47348
rect 27636 47292 34300 47348
rect 34356 47292 34366 47348
rect 20132 47236 20188 47292
rect 8530 47180 8540 47236
rect 8596 47180 10556 47236
rect 10612 47180 10622 47236
rect 12338 47180 12348 47236
rect 12404 47180 15820 47236
rect 15876 47180 15886 47236
rect 16034 47180 16044 47236
rect 16100 47180 19012 47236
rect 20132 47180 29148 47236
rect 29204 47180 29214 47236
rect 30370 47180 30380 47236
rect 30436 47180 30828 47236
rect 30884 47180 30894 47236
rect 31938 47180 31948 47236
rect 32004 47180 33068 47236
rect 33124 47180 33134 47236
rect 33282 47180 33292 47236
rect 33348 47180 38668 47236
rect 18956 47124 19012 47180
rect 38612 47124 38668 47180
rect 2146 47068 2156 47124
rect 2212 47068 4956 47124
rect 5012 47068 5022 47124
rect 6514 47068 6524 47124
rect 6580 47068 8316 47124
rect 8372 47068 8382 47124
rect 8530 47068 8540 47124
rect 8596 47068 10164 47124
rect 10322 47068 10332 47124
rect 10388 47068 18732 47124
rect 18788 47068 18798 47124
rect 18956 47068 24052 47124
rect 24210 47068 24220 47124
rect 24276 47068 27468 47124
rect 27524 47068 27534 47124
rect 27794 47068 27804 47124
rect 27860 47068 36204 47124
rect 36260 47068 36270 47124
rect 38612 47068 40348 47124
rect 40404 47068 40414 47124
rect 10108 47012 10164 47068
rect 23996 47012 24052 47068
rect 8306 46956 8316 47012
rect 8372 46844 8428 47012
rect 10108 46956 12124 47012
rect 12180 46956 12190 47012
rect 23996 46956 24556 47012
rect 24612 46956 24622 47012
rect 8484 46844 8494 46900
rect 12674 46844 12684 46900
rect 12740 46844 27020 46900
rect 27076 46844 27086 46900
rect 8306 46732 8316 46788
rect 8372 46732 19852 46788
rect 19908 46732 19918 46788
rect 7186 46620 7196 46676
rect 7252 46620 15260 46676
rect 15316 46620 15326 46676
rect 17938 46620 17948 46676
rect 18004 46620 29932 46676
rect 29988 46620 29998 46676
rect 27570 46508 27580 46564
rect 27636 46508 29260 46564
rect 29316 46508 32284 46564
rect 32340 46508 38668 46564
rect 38612 46452 38668 46508
rect 5842 46396 5852 46452
rect 5908 46396 10780 46452
rect 10836 46396 10846 46452
rect 12226 46396 12236 46452
rect 12292 46396 13356 46452
rect 13412 46396 13422 46452
rect 27682 46396 27692 46452
rect 27748 46396 37548 46452
rect 37604 46396 37614 46452
rect 38612 46396 39340 46452
rect 39396 46396 39406 46452
rect 49200 46368 49800 46480
rect 10322 46284 10332 46340
rect 10388 46284 12796 46340
rect 12852 46284 12862 46340
rect 13020 46284 22204 46340
rect 22260 46284 22270 46340
rect 30594 46284 30604 46340
rect 30660 46284 31052 46340
rect 31108 46284 31118 46340
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 13020 46228 13076 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 9762 46172 9772 46228
rect 9828 46172 13076 46228
rect 13346 46172 13356 46228
rect 13412 46172 28364 46228
rect 28420 46172 33628 46228
rect 33684 46172 33694 46228
rect 11666 46060 11676 46116
rect 11732 46060 11788 46116
rect 11844 46060 11854 46116
rect 13234 46060 13244 46116
rect 13300 46060 27692 46116
rect 27748 46060 27758 46116
rect 28018 46060 28028 46116
rect 28084 46060 33628 46116
rect 33684 46060 33694 46116
rect 7298 45948 7308 46004
rect 7364 45948 17388 46004
rect 17444 45948 17454 46004
rect 17686 45948 17724 46004
rect 17780 45948 17790 46004
rect 22866 45948 22876 46004
rect 22932 45948 27692 46004
rect 27748 45948 27758 46004
rect 27906 45948 27916 46004
rect 27972 45948 33852 46004
rect 33908 45948 33918 46004
rect 10882 45836 10892 45892
rect 10948 45836 11452 45892
rect 11508 45836 13580 45892
rect 13636 45836 13646 45892
rect 16594 45836 16604 45892
rect 16660 45836 20188 45892
rect 24546 45836 24556 45892
rect 24612 45836 27356 45892
rect 27412 45836 32172 45892
rect 32228 45836 32238 45892
rect 35858 45836 35868 45892
rect 35924 45836 36092 45892
rect 36148 45836 41804 45892
rect 41860 45836 41870 45892
rect 200 45780 800 45808
rect 20132 45780 20188 45836
rect 200 45724 1708 45780
rect 1764 45724 1774 45780
rect 2594 45724 2604 45780
rect 2660 45724 10836 45780
rect 10994 45724 11004 45780
rect 11060 45724 18172 45780
rect 18228 45724 18238 45780
rect 20132 45724 25676 45780
rect 25732 45724 25742 45780
rect 26898 45724 26908 45780
rect 26964 45724 30156 45780
rect 30212 45724 30222 45780
rect 30930 45724 30940 45780
rect 30996 45724 31500 45780
rect 31556 45724 41356 45780
rect 41412 45724 41422 45780
rect 200 45696 800 45724
rect 10780 45668 10836 45724
rect 8194 45612 8204 45668
rect 8260 45612 8540 45668
rect 8596 45612 8606 45668
rect 10780 45612 11508 45668
rect 11778 45612 11788 45668
rect 11844 45612 12348 45668
rect 12404 45612 12414 45668
rect 13458 45612 13468 45668
rect 13524 45612 20916 45668
rect 27682 45612 27692 45668
rect 27748 45612 28364 45668
rect 28420 45612 28430 45668
rect 29586 45612 29596 45668
rect 29652 45612 31500 45668
rect 31556 45612 31566 45668
rect 32162 45612 32172 45668
rect 32228 45612 37100 45668
rect 37156 45612 40572 45668
rect 40628 45612 40638 45668
rect 40898 45612 40908 45668
rect 40964 45612 47740 45668
rect 47796 45612 47806 45668
rect 4284 45500 11228 45556
rect 11284 45500 11294 45556
rect 4284 45332 4340 45500
rect 11452 45444 11508 45612
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 20860 45444 20916 45612
rect 27794 45500 27804 45556
rect 27860 45500 28028 45556
rect 28084 45500 28094 45556
rect 29250 45500 29260 45556
rect 29316 45500 29484 45556
rect 29540 45500 29550 45556
rect 29782 45500 29820 45556
rect 29876 45500 29886 45556
rect 30146 45500 30156 45556
rect 30212 45500 35644 45556
rect 35700 45500 35710 45556
rect 11442 45388 11452 45444
rect 11508 45388 12460 45444
rect 12516 45388 12526 45444
rect 15250 45388 15260 45444
rect 15316 45388 16604 45444
rect 16660 45388 16670 45444
rect 20850 45388 20860 45444
rect 20916 45388 27132 45444
rect 27188 45388 27198 45444
rect 27458 45388 27468 45444
rect 27524 45388 28700 45444
rect 28756 45388 28766 45444
rect 30258 45388 30268 45444
rect 30324 45388 37212 45444
rect 37268 45388 37278 45444
rect 4274 45276 4284 45332
rect 4340 45276 4350 45332
rect 4610 45276 4620 45332
rect 4676 45276 13244 45332
rect 13300 45276 15148 45332
rect 15204 45276 15214 45332
rect 19506 45276 19516 45332
rect 19572 45276 20636 45332
rect 20692 45276 21532 45332
rect 21588 45276 21598 45332
rect 27010 45276 27020 45332
rect 27076 45276 31500 45332
rect 31556 45276 31566 45332
rect 7830 45164 7868 45220
rect 7924 45164 7934 45220
rect 10098 45164 10108 45220
rect 10164 45164 11116 45220
rect 11172 45164 14700 45220
rect 14756 45164 14766 45220
rect 18610 45164 18620 45220
rect 18676 45164 20188 45220
rect 20244 45164 20254 45220
rect 22978 45164 22988 45220
rect 23044 45164 24892 45220
rect 24948 45164 24958 45220
rect 28018 45164 28028 45220
rect 28084 45164 34860 45220
rect 34916 45164 34926 45220
rect 6290 45052 6300 45108
rect 6356 45052 6748 45108
rect 6804 45052 6814 45108
rect 7942 45052 7980 45108
rect 8036 45052 8046 45108
rect 9874 45052 9884 45108
rect 9940 45052 11172 45108
rect 11330 45052 11340 45108
rect 11396 45052 11452 45108
rect 11508 45052 11518 45108
rect 11666 45052 11676 45108
rect 11732 45052 11788 45108
rect 11844 45052 11854 45108
rect 14018 45052 14028 45108
rect 14084 45052 15372 45108
rect 15428 45052 15438 45108
rect 16706 45052 16716 45108
rect 16772 45052 17724 45108
rect 17780 45052 17790 45108
rect 19590 45052 19628 45108
rect 19684 45052 19694 45108
rect 28102 45052 28140 45108
rect 28196 45052 28206 45108
rect 29698 45052 29708 45108
rect 29764 45052 30044 45108
rect 30100 45052 30110 45108
rect 30818 45052 30828 45108
rect 30884 45052 33404 45108
rect 33460 45052 33470 45108
rect 33618 45052 33628 45108
rect 33684 45052 38220 45108
rect 38276 45052 38286 45108
rect 11116 44996 11172 45052
rect 49200 45024 49800 45136
rect 1922 44940 1932 44996
rect 1988 44940 10892 44996
rect 10948 44940 10958 44996
rect 11116 44940 12908 44996
rect 12964 44940 14756 44996
rect 18834 44940 18844 44996
rect 18900 44940 27580 44996
rect 27636 44940 27646 44996
rect 28354 44940 28364 44996
rect 28420 44940 29708 44996
rect 29764 44940 29774 44996
rect 30146 44940 30156 44996
rect 30212 44940 31052 44996
rect 31108 44940 31118 44996
rect 36866 44940 36876 44996
rect 36932 44940 37548 44996
rect 37604 44940 37614 44996
rect 14700 44884 14756 44940
rect 3714 44828 3724 44884
rect 3780 44828 10556 44884
rect 10612 44828 11452 44884
rect 11508 44828 11518 44884
rect 12310 44828 12348 44884
rect 12404 44828 12414 44884
rect 13458 44828 13468 44884
rect 13524 44828 14644 44884
rect 14700 44828 21868 44884
rect 21924 44828 21934 44884
rect 22642 44828 22652 44884
rect 22708 44828 29372 44884
rect 29428 44828 37772 44884
rect 37828 44828 38332 44884
rect 38388 44828 38398 44884
rect 14588 44772 14644 44828
rect 9762 44716 9772 44772
rect 9828 44716 14364 44772
rect 14420 44716 14430 44772
rect 14588 44716 22428 44772
rect 22484 44716 24780 44772
rect 24836 44716 24846 44772
rect 24994 44716 25004 44772
rect 25060 44716 26684 44772
rect 26740 44716 28308 44772
rect 29474 44716 29484 44772
rect 29540 44716 31052 44772
rect 31108 44716 34020 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 28252 44660 28308 44716
rect 5506 44604 5516 44660
rect 5572 44604 12348 44660
rect 12404 44604 12414 44660
rect 14018 44604 14028 44660
rect 14084 44604 21196 44660
rect 21252 44604 28028 44660
rect 28084 44604 28094 44660
rect 28252 44604 30268 44660
rect 30324 44604 30334 44660
rect 30930 44604 30940 44660
rect 30996 44604 33740 44660
rect 33796 44604 33806 44660
rect 33964 44548 34020 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 7298 44492 7308 44548
rect 7364 44492 9772 44548
rect 9828 44492 9838 44548
rect 10210 44492 10220 44548
rect 10276 44492 20412 44548
rect 20468 44492 20478 44548
rect 31154 44492 31164 44548
rect 31220 44492 31388 44548
rect 31444 44492 31454 44548
rect 31602 44492 31612 44548
rect 31668 44492 31836 44548
rect 31892 44492 31902 44548
rect 33964 44492 35308 44548
rect 35364 44492 35374 44548
rect 4134 44380 4172 44436
rect 4228 44380 4238 44436
rect 6738 44380 6748 44436
rect 6804 44380 14812 44436
rect 14868 44380 14878 44436
rect 22194 44380 22204 44436
rect 22260 44380 24556 44436
rect 24612 44380 25340 44436
rect 25396 44380 25406 44436
rect 25890 44380 25900 44436
rect 25956 44380 35532 44436
rect 35588 44380 35598 44436
rect 35746 44380 35756 44436
rect 35812 44380 40460 44436
rect 40516 44380 40526 44436
rect 4610 44268 4620 44324
rect 4676 44268 11564 44324
rect 11620 44268 12908 44324
rect 12964 44268 12974 44324
rect 13132 44268 14700 44324
rect 14756 44268 14766 44324
rect 15362 44268 15372 44324
rect 15428 44268 17724 44324
rect 17780 44268 17948 44324
rect 18004 44268 19516 44324
rect 19572 44268 19582 44324
rect 28690 44268 28700 44324
rect 28756 44268 29484 44324
rect 29540 44268 29550 44324
rect 29698 44268 29708 44324
rect 29764 44268 38780 44324
rect 38836 44268 38846 44324
rect 13132 44212 13188 44268
rect 4274 44156 4284 44212
rect 4340 44156 4956 44212
rect 5012 44156 5022 44212
rect 5842 44156 5852 44212
rect 5908 44156 10332 44212
rect 10388 44156 10398 44212
rect 10556 44156 13188 44212
rect 13794 44156 13804 44212
rect 13860 44156 16044 44212
rect 16100 44156 16110 44212
rect 25106 44156 25116 44212
rect 25172 44156 28364 44212
rect 28420 44156 28430 44212
rect 28802 44156 28812 44212
rect 28868 44156 32788 44212
rect 35298 44156 35308 44212
rect 35364 44156 38332 44212
rect 38388 44156 38398 44212
rect 10556 44100 10612 44156
rect 32732 44100 32788 44156
rect 38612 44100 38668 44212
rect 38724 44156 38734 44212
rect 6290 44044 6300 44100
rect 6356 44044 8428 44100
rect 8484 44044 8494 44100
rect 8950 44044 8988 44100
rect 9044 44044 9054 44100
rect 10332 44044 10612 44100
rect 10770 44044 10780 44100
rect 10836 44044 12572 44100
rect 12628 44044 18844 44100
rect 18900 44044 18910 44100
rect 19068 44044 23660 44100
rect 23716 44044 23726 44100
rect 26684 44044 27692 44100
rect 27748 44044 29708 44100
rect 29764 44044 29774 44100
rect 30034 44044 30044 44100
rect 30100 44044 31724 44100
rect 31780 44044 31790 44100
rect 32722 44044 32732 44100
rect 32788 44044 34524 44100
rect 34580 44044 36652 44100
rect 36708 44044 36718 44100
rect 38444 44044 38668 44100
rect 10332 43876 10388 44044
rect 19068 43988 19124 44044
rect 26684 43988 26740 44044
rect 38444 43988 38500 44044
rect 10546 43932 10556 43988
rect 10612 43932 11396 43988
rect 11778 43932 11788 43988
rect 11844 43932 12124 43988
rect 12180 43932 14980 43988
rect 15698 43932 15708 43988
rect 15764 43932 19124 43988
rect 22530 43932 22540 43988
rect 22596 43932 26740 43988
rect 26852 43932 30380 43988
rect 30436 43932 34412 43988
rect 34468 43932 34972 43988
rect 35028 43932 35038 43988
rect 36652 43932 38500 43988
rect 7634 43820 7644 43876
rect 7700 43820 10388 43876
rect 200 43764 800 43792
rect 11340 43764 11396 43932
rect 14924 43876 14980 43932
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 26852 43876 26908 43932
rect 36652 43876 36708 43932
rect 14924 43820 18956 43876
rect 19012 43820 19022 43876
rect 20178 43820 20188 43876
rect 20244 43820 26908 43876
rect 29362 43820 29372 43876
rect 29428 43820 29484 43876
rect 29540 43820 34412 43876
rect 34468 43820 34478 43876
rect 34850 43820 34860 43876
rect 34916 43820 36708 43876
rect 36866 43820 36876 43876
rect 36932 43820 37884 43876
rect 37940 43820 39900 43876
rect 39956 43820 39966 43876
rect 200 43708 2156 43764
rect 2212 43708 2222 43764
rect 10630 43708 10668 43764
rect 10724 43708 10734 43764
rect 11330 43708 11340 43764
rect 11396 43708 11406 43764
rect 11554 43708 11564 43764
rect 11620 43708 11900 43764
rect 11956 43708 11966 43764
rect 12338 43708 12348 43764
rect 12404 43708 12460 43764
rect 12516 43708 12526 43764
rect 15138 43708 15148 43764
rect 15204 43708 25900 43764
rect 25956 43708 25966 43764
rect 27682 43708 27692 43764
rect 27748 43708 29036 43764
rect 29092 43708 29102 43764
rect 30482 43708 30492 43764
rect 30548 43708 32396 43764
rect 32452 43708 32462 43764
rect 33506 43708 33516 43764
rect 33572 43708 38108 43764
rect 38164 43708 38174 43764
rect 38322 43708 38332 43764
rect 38388 43708 38892 43764
rect 38948 43708 38958 43764
rect 200 43680 800 43708
rect 4946 43596 4956 43652
rect 5012 43596 6300 43652
rect 6356 43596 6636 43652
rect 6692 43596 6702 43652
rect 6850 43596 6860 43652
rect 6916 43596 8204 43652
rect 8260 43596 8270 43652
rect 10770 43596 10780 43652
rect 10836 43596 11788 43652
rect 11844 43596 11854 43652
rect 13682 43596 13692 43652
rect 13748 43596 14588 43652
rect 14644 43596 14654 43652
rect 14802 43596 14812 43652
rect 14868 43596 14906 43652
rect 17826 43596 17836 43652
rect 17892 43596 18396 43652
rect 18452 43596 18462 43652
rect 22194 43596 22204 43652
rect 22260 43596 22652 43652
rect 22708 43596 22718 43652
rect 30034 43596 30044 43652
rect 30100 43596 30268 43652
rect 30324 43596 30334 43652
rect 30528 43596 30604 43652
rect 30660 43596 35756 43652
rect 35812 43596 35822 43652
rect 36754 43596 36764 43652
rect 36820 43596 39228 43652
rect 39284 43596 39294 43652
rect 4162 43484 4172 43540
rect 4228 43484 11228 43540
rect 11284 43484 11294 43540
rect 11666 43484 11676 43540
rect 11732 43484 12460 43540
rect 12516 43484 12526 43540
rect 14018 43484 14028 43540
rect 14084 43484 14476 43540
rect 14532 43484 14542 43540
rect 17042 43484 17052 43540
rect 17108 43484 20188 43540
rect 24070 43484 24108 43540
rect 24164 43484 24174 43540
rect 24546 43484 24556 43540
rect 24612 43484 30940 43540
rect 30996 43484 31006 43540
rect 31238 43484 31276 43540
rect 31332 43484 31342 43540
rect 31490 43484 31500 43540
rect 31556 43484 31836 43540
rect 31892 43484 31902 43540
rect 32498 43484 32508 43540
rect 32564 43484 33684 43540
rect 34738 43484 34748 43540
rect 34804 43484 35756 43540
rect 35812 43484 35822 43540
rect 37986 43484 37996 43540
rect 38052 43484 39676 43540
rect 39732 43484 39742 43540
rect 20132 43428 20188 43484
rect 33628 43428 33684 43484
rect 2706 43372 2716 43428
rect 2772 43372 8652 43428
rect 8708 43372 10668 43428
rect 10724 43372 10734 43428
rect 13692 43372 17276 43428
rect 17332 43372 17612 43428
rect 17668 43372 17678 43428
rect 17938 43372 17948 43428
rect 18004 43372 18060 43428
rect 18116 43372 18126 43428
rect 20132 43372 21532 43428
rect 21588 43372 21598 43428
rect 23538 43372 23548 43428
rect 23604 43372 24444 43428
rect 24500 43372 24510 43428
rect 28998 43372 29036 43428
rect 29092 43372 29102 43428
rect 29810 43372 29820 43428
rect 29876 43372 30212 43428
rect 30370 43372 30380 43428
rect 30436 43372 33068 43428
rect 33124 43372 33134 43428
rect 33628 43372 39788 43428
rect 39844 43372 39854 43428
rect 13692 43316 13748 43372
rect 30156 43316 30212 43372
rect 3378 43260 3388 43316
rect 3444 43260 4620 43316
rect 4676 43260 5348 43316
rect 5506 43260 5516 43316
rect 5572 43260 13692 43316
rect 13748 43260 13758 43316
rect 16930 43260 16940 43316
rect 16996 43260 27804 43316
rect 27860 43260 27870 43316
rect 28914 43260 28924 43316
rect 28980 43260 29708 43316
rect 29764 43260 29774 43316
rect 29894 43260 29932 43316
rect 29988 43260 29998 43316
rect 30156 43260 34188 43316
rect 34244 43260 36652 43316
rect 36708 43260 36718 43316
rect 37426 43260 37436 43316
rect 37492 43260 37548 43316
rect 37604 43260 40348 43316
rect 40404 43260 40414 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 5292 43092 5348 43260
rect 7298 43148 7308 43204
rect 7364 43148 14196 43204
rect 17378 43148 17388 43204
rect 17444 43148 19404 43204
rect 19460 43148 19470 43204
rect 22642 43148 22652 43204
rect 22708 43148 31836 43204
rect 31892 43148 31902 43204
rect 32386 43148 32396 43204
rect 32452 43148 33516 43204
rect 33572 43148 33582 43204
rect 33730 43148 33740 43204
rect 33796 43148 34748 43204
rect 34804 43148 34814 43204
rect 35746 43148 35756 43204
rect 35812 43148 36876 43204
rect 36932 43148 36942 43204
rect 5292 43036 12684 43092
rect 12740 43036 12750 43092
rect 14140 42980 14196 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 49200 43092 49800 43120
rect 14354 43036 14364 43092
rect 14420 43036 21980 43092
rect 22036 43036 23772 43092
rect 23828 43036 23838 43092
rect 26898 43036 26908 43092
rect 26964 43036 34076 43092
rect 34132 43036 34860 43092
rect 34916 43036 34926 43092
rect 36166 43036 36204 43092
rect 36260 43036 36270 43092
rect 47282 43036 47292 43092
rect 47348 43036 48076 43092
rect 48132 43036 49800 43092
rect 34860 42980 34916 43036
rect 49200 43008 49800 43036
rect 4050 42924 4060 42980
rect 4116 42924 7084 42980
rect 7140 42924 8428 42980
rect 14140 42924 18060 42980
rect 18116 42924 18126 42980
rect 25330 42924 25340 42980
rect 25396 42924 32732 42980
rect 32788 42924 32798 42980
rect 33506 42924 33516 42980
rect 33572 42924 34524 42980
rect 34580 42924 34590 42980
rect 34860 42924 35532 42980
rect 35588 42924 35598 42980
rect 8372 42868 8428 42924
rect 2818 42812 2828 42868
rect 2884 42812 6524 42868
rect 6580 42812 6590 42868
rect 8372 42812 9996 42868
rect 10052 42812 12012 42868
rect 12068 42812 15036 42868
rect 15092 42812 15102 42868
rect 17378 42812 17388 42868
rect 17444 42812 20188 42868
rect 20244 42812 20254 42868
rect 20402 42812 20412 42868
rect 20468 42812 20860 42868
rect 20916 42812 20972 42868
rect 21028 42812 21038 42868
rect 28578 42812 28588 42868
rect 28644 42812 29372 42868
rect 29428 42812 29438 42868
rect 29810 42812 29820 42868
rect 29876 42812 30156 42868
rect 30212 42812 35252 42868
rect 35308 42812 35318 42868
rect 39330 42812 39340 42868
rect 39396 42812 40124 42868
rect 40180 42812 40190 42868
rect 4162 42700 4172 42756
rect 4228 42700 9884 42756
rect 9940 42700 9950 42756
rect 18946 42700 18956 42756
rect 19012 42700 21644 42756
rect 21700 42700 21710 42756
rect 24546 42700 24556 42756
rect 24612 42700 25116 42756
rect 25172 42700 25182 42756
rect 27906 42700 27916 42756
rect 27972 42700 28476 42756
rect 28532 42700 28542 42756
rect 28914 42700 28924 42756
rect 28980 42700 29708 42756
rect 29764 42700 30380 42756
rect 30436 42700 30446 42756
rect 31154 42700 31164 42756
rect 31220 42700 31276 42756
rect 31332 42700 31342 42756
rect 31490 42700 31500 42756
rect 31556 42700 35308 42756
rect 35634 42700 35644 42756
rect 35700 42700 36652 42756
rect 36708 42700 36718 42756
rect 35252 42644 35308 42700
rect 8166 42588 8204 42644
rect 8260 42588 8270 42644
rect 9062 42588 9100 42644
rect 9156 42588 9166 42644
rect 11442 42588 11452 42644
rect 11508 42588 17052 42644
rect 17108 42588 17118 42644
rect 23762 42588 23772 42644
rect 23828 42588 30604 42644
rect 30660 42588 30670 42644
rect 30930 42588 30940 42644
rect 30996 42588 31388 42644
rect 31444 42588 31454 42644
rect 31602 42588 31612 42644
rect 31668 42588 31706 42644
rect 31826 42588 31836 42644
rect 31892 42588 33068 42644
rect 33124 42588 33134 42644
rect 33282 42588 33292 42644
rect 33348 42588 34972 42644
rect 35028 42588 35038 42644
rect 35252 42588 37436 42644
rect 37492 42588 37502 42644
rect 37660 42588 40124 42644
rect 40180 42588 40190 42644
rect 37660 42532 37716 42588
rect 3714 42476 3724 42532
rect 3780 42476 8764 42532
rect 8820 42476 8988 42532
rect 9044 42476 9054 42532
rect 9286 42476 9324 42532
rect 9380 42476 9390 42532
rect 10434 42476 10444 42532
rect 10500 42476 23548 42532
rect 23604 42476 23614 42532
rect 25218 42476 25228 42532
rect 25284 42476 29820 42532
rect 29876 42476 29886 42532
rect 30370 42476 30380 42532
rect 30436 42476 32340 42532
rect 32498 42476 32508 42532
rect 32564 42476 32956 42532
rect 33012 42476 33022 42532
rect 33954 42476 33964 42532
rect 34020 42476 34860 42532
rect 34916 42476 37716 42532
rect 38098 42476 38108 42532
rect 38164 42476 38668 42532
rect 38724 42476 38734 42532
rect 39218 42476 39228 42532
rect 39284 42476 39452 42532
rect 39508 42476 39518 42532
rect 200 42420 800 42448
rect 200 42364 1820 42420
rect 1876 42364 1886 42420
rect 4610 42364 4620 42420
rect 4676 42364 13916 42420
rect 13972 42364 13982 42420
rect 14690 42364 14700 42420
rect 14756 42364 14812 42420
rect 14868 42364 18508 42420
rect 18564 42364 18574 42420
rect 20850 42364 20860 42420
rect 20916 42364 25788 42420
rect 25844 42364 25854 42420
rect 29026 42364 29036 42420
rect 29092 42364 30716 42420
rect 30772 42364 30782 42420
rect 200 42336 800 42364
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 32284 42308 32340 42476
rect 33394 42364 33404 42420
rect 33460 42364 34972 42420
rect 35028 42364 35038 42420
rect 35746 42364 35756 42420
rect 35812 42364 40572 42420
rect 40628 42364 40638 42420
rect 9762 42252 9772 42308
rect 9828 42252 9996 42308
rect 10052 42252 10062 42308
rect 10546 42252 10556 42308
rect 10612 42252 12796 42308
rect 12852 42252 12862 42308
rect 13356 42252 18956 42308
rect 19012 42252 19022 42308
rect 21186 42252 21196 42308
rect 21252 42252 26124 42308
rect 26180 42252 28588 42308
rect 28644 42252 28654 42308
rect 31500 42252 31948 42308
rect 32004 42252 32014 42308
rect 32284 42252 36204 42308
rect 36260 42252 36270 42308
rect 2706 42140 2716 42196
rect 2772 42140 3164 42196
rect 3220 42140 3230 42196
rect 3612 42140 7868 42196
rect 7924 42140 10444 42196
rect 10500 42140 10510 42196
rect 10658 42140 10668 42196
rect 10724 42140 12124 42196
rect 12180 42140 12190 42196
rect 3612 42084 3668 42140
rect 2370 42028 2380 42084
rect 2436 42028 3612 42084
rect 3668 42028 3678 42084
rect 6934 42028 6972 42084
rect 7028 42028 7038 42084
rect 8530 42028 8540 42084
rect 8596 42028 9212 42084
rect 9268 42028 9278 42084
rect 9874 42028 9884 42084
rect 9940 42028 10892 42084
rect 10948 42028 10958 42084
rect 13356 41972 13412 42252
rect 18050 42140 18060 42196
rect 18116 42140 18172 42196
rect 18228 42140 18238 42196
rect 18386 42140 18396 42196
rect 18452 42140 24948 42196
rect 25106 42140 25116 42196
rect 25172 42140 25788 42196
rect 25844 42140 26908 42196
rect 26964 42140 26974 42196
rect 28690 42140 28700 42196
rect 28756 42140 31164 42196
rect 31220 42140 31230 42196
rect 24892 42084 24948 42140
rect 14578 42028 14588 42084
rect 14644 42028 15596 42084
rect 15652 42028 15662 42084
rect 16930 42028 16940 42084
rect 16996 42028 17836 42084
rect 17892 42028 18732 42084
rect 18788 42028 18798 42084
rect 19058 42028 19068 42084
rect 19124 42028 22876 42084
rect 22932 42028 22942 42084
rect 23090 42028 23100 42084
rect 23156 42028 23884 42084
rect 23940 42028 24500 42084
rect 24892 42028 28700 42084
rect 28756 42028 29036 42084
rect 29092 42028 29484 42084
rect 29540 42028 29550 42084
rect 29922 42028 29932 42084
rect 29988 42028 31276 42084
rect 31332 42028 31342 42084
rect 24444 41972 24500 42028
rect 31500 41972 31556 42252
rect 32834 42140 32844 42196
rect 32900 42140 33068 42196
rect 33124 42140 33134 42196
rect 33404 42140 35476 42196
rect 33404 42084 33460 42140
rect 35420 42084 35476 42140
rect 31910 42028 31948 42084
rect 32004 42028 32014 42084
rect 32162 42028 32172 42084
rect 32228 42028 33460 42084
rect 34710 42028 34748 42084
rect 34804 42028 34814 42084
rect 35420 42028 37044 42084
rect 38434 42028 38444 42084
rect 38500 42028 39004 42084
rect 39060 42028 39070 42084
rect 36988 41972 37044 42028
rect 2146 41916 2156 41972
rect 2212 41916 6188 41972
rect 6244 41916 6254 41972
rect 6402 41916 6412 41972
rect 6468 41916 6636 41972
rect 6692 41916 6702 41972
rect 6850 41916 6860 41972
rect 6916 41916 7756 41972
rect 7812 41916 7822 41972
rect 8754 41916 8764 41972
rect 8820 41916 13412 41972
rect 18162 41916 18172 41972
rect 18228 41916 18396 41972
rect 18452 41916 19516 41972
rect 19572 41916 19582 41972
rect 22082 41916 22092 41972
rect 22148 41916 22316 41972
rect 22372 41916 22382 41972
rect 24434 41916 24444 41972
rect 24500 41916 24510 41972
rect 26898 41916 26908 41972
rect 26964 41916 29484 41972
rect 29540 41916 29550 41972
rect 29782 41916 29820 41972
rect 29876 41916 29886 41972
rect 30034 41916 30044 41972
rect 30100 41916 30716 41972
rect 30772 41916 31556 41972
rect 31826 41916 31836 41972
rect 31892 41916 35308 41972
rect 35364 41916 35644 41972
rect 35700 41916 35710 41972
rect 35970 41916 35980 41972
rect 36036 41916 36764 41972
rect 36820 41916 36830 41972
rect 36978 41916 36988 41972
rect 37044 41916 38668 41972
rect 38612 41860 38668 41916
rect 3462 41804 3500 41860
rect 3556 41804 3566 41860
rect 4386 41804 4396 41860
rect 4452 41804 4956 41860
rect 5012 41804 5022 41860
rect 5180 41804 8316 41860
rect 8372 41804 8382 41860
rect 8866 41804 8876 41860
rect 8932 41804 9548 41860
rect 9604 41804 9614 41860
rect 9762 41804 9772 41860
rect 9828 41804 16716 41860
rect 16772 41804 19964 41860
rect 20020 41804 20030 41860
rect 20132 41804 23324 41860
rect 23380 41804 23390 41860
rect 23538 41804 23548 41860
rect 23604 41804 31164 41860
rect 31220 41804 32172 41860
rect 32228 41804 32238 41860
rect 32610 41804 32620 41860
rect 32676 41804 37436 41860
rect 37492 41804 37502 41860
rect 38612 41804 39116 41860
rect 39172 41804 39182 41860
rect 5180 41748 5236 41804
rect 20132 41748 20188 41804
rect 2818 41692 2828 41748
rect 2884 41692 5236 41748
rect 5954 41692 5964 41748
rect 6020 41692 6636 41748
rect 6692 41692 6702 41748
rect 7298 41692 7308 41748
rect 7364 41692 9884 41748
rect 9940 41692 9950 41748
rect 13122 41692 13132 41748
rect 13188 41692 13468 41748
rect 13524 41692 13534 41748
rect 19506 41692 19516 41748
rect 19572 41692 20188 41748
rect 21410 41692 21420 41748
rect 21476 41692 22092 41748
rect 22148 41692 22158 41748
rect 30342 41692 30380 41748
rect 30436 41692 30446 41748
rect 31378 41692 31388 41748
rect 31444 41692 33292 41748
rect 33348 41692 33358 41748
rect 33506 41692 33516 41748
rect 33572 41692 33610 41748
rect 34962 41692 34972 41748
rect 35028 41692 35084 41748
rect 35140 41692 40460 41748
rect 40516 41692 40526 41748
rect 4834 41580 4844 41636
rect 4900 41580 9436 41636
rect 9492 41580 9502 41636
rect 10770 41580 10780 41636
rect 10836 41580 27356 41636
rect 27412 41580 27422 41636
rect 28578 41580 28588 41636
rect 28644 41580 32060 41636
rect 32116 41580 32126 41636
rect 32498 41580 32508 41636
rect 32564 41580 33404 41636
rect 33460 41580 33470 41636
rect 34066 41580 34076 41636
rect 34132 41580 34636 41636
rect 34692 41580 34702 41636
rect 35634 41580 35644 41636
rect 35700 41580 42028 41636
rect 42084 41580 42094 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 3266 41468 3276 41524
rect 3332 41468 4116 41524
rect 6626 41468 6636 41524
rect 6692 41468 11340 41524
rect 11396 41468 11406 41524
rect 12114 41468 12124 41524
rect 12180 41468 17052 41524
rect 17108 41468 19180 41524
rect 19236 41468 20188 41524
rect 4060 41412 4116 41468
rect 20132 41412 20188 41468
rect 26852 41468 28812 41524
rect 28868 41468 29148 41524
rect 29204 41468 29214 41524
rect 30034 41468 30044 41524
rect 30100 41468 30156 41524
rect 30212 41468 34188 41524
rect 34244 41468 34254 41524
rect 35634 41468 35644 41524
rect 35700 41468 35868 41524
rect 35924 41468 35934 41524
rect 26852 41412 26908 41468
rect 4050 41356 4060 41412
rect 4116 41356 5628 41412
rect 5684 41356 7980 41412
rect 8036 41356 8046 41412
rect 8614 41356 8652 41412
rect 8708 41356 8718 41412
rect 8866 41356 8876 41412
rect 8932 41356 15260 41412
rect 15316 41356 15820 41412
rect 15876 41356 15886 41412
rect 20132 41356 20972 41412
rect 21028 41356 21038 41412
rect 24994 41356 25004 41412
rect 25060 41356 26908 41412
rect 28242 41356 28252 41412
rect 28308 41356 33180 41412
rect 33236 41356 33246 41412
rect 34626 41356 34636 41412
rect 34692 41356 40572 41412
rect 40628 41356 40638 41412
rect 3938 41244 3948 41300
rect 4004 41244 5964 41300
rect 6020 41244 8988 41300
rect 9044 41244 9054 41300
rect 9314 41244 9324 41300
rect 9380 41244 9548 41300
rect 9604 41244 9614 41300
rect 10546 41244 10556 41300
rect 10612 41244 12908 41300
rect 12964 41244 14140 41300
rect 14196 41244 14206 41300
rect 14466 41244 14476 41300
rect 14532 41244 15148 41300
rect 15204 41244 15214 41300
rect 17378 41244 17388 41300
rect 17444 41244 24052 41300
rect 24210 41244 24220 41300
rect 24276 41244 26908 41300
rect 26964 41244 26974 41300
rect 29250 41244 29260 41300
rect 29316 41244 29372 41300
rect 29428 41244 29438 41300
rect 29558 41244 29596 41300
rect 29652 41244 29662 41300
rect 30818 41244 30828 41300
rect 30884 41244 31500 41300
rect 31556 41244 31566 41300
rect 31826 41244 31836 41300
rect 31892 41244 34412 41300
rect 34468 41244 35196 41300
rect 35252 41244 35262 41300
rect 35634 41244 35644 41300
rect 35700 41244 36092 41300
rect 36148 41244 36158 41300
rect 23996 41188 24052 41244
rect 2370 41132 2380 41188
rect 2436 41132 8036 41188
rect 8306 41132 8316 41188
rect 8372 41132 8652 41188
rect 8708 41132 8718 41188
rect 9090 41132 9100 41188
rect 9156 41132 9166 41188
rect 9650 41132 9660 41188
rect 9716 41132 14588 41188
rect 14644 41132 14654 41188
rect 16482 41132 16492 41188
rect 16548 41132 17500 41188
rect 17556 41132 17566 41188
rect 19954 41132 19964 41188
rect 20020 41132 21196 41188
rect 21252 41132 21262 41188
rect 23538 41132 23548 41188
rect 23604 41132 23660 41188
rect 23716 41132 23726 41188
rect 23996 41132 26460 41188
rect 26516 41132 26526 41188
rect 27906 41132 27916 41188
rect 27972 41132 32396 41188
rect 32452 41132 32462 41188
rect 32610 41132 32620 41188
rect 32676 41132 33068 41188
rect 33124 41132 33134 41188
rect 33328 41132 33404 41188
rect 33460 41132 34804 41188
rect 34962 41132 34972 41188
rect 35028 41132 36652 41188
rect 36708 41132 36718 41188
rect 7980 41076 8036 41132
rect 9100 41076 9156 41132
rect 34748 41076 34804 41132
rect 3490 41020 3500 41076
rect 3556 41020 4844 41076
rect 4900 41020 4910 41076
rect 6962 41020 6972 41076
rect 7028 41020 7308 41076
rect 7364 41020 7374 41076
rect 7980 41020 9156 41076
rect 9212 41020 9996 41076
rect 10052 41020 14028 41076
rect 14084 41020 14094 41076
rect 17266 41020 17276 41076
rect 17332 41020 18172 41076
rect 18228 41020 18238 41076
rect 20178 41020 20188 41076
rect 20244 41020 20860 41076
rect 20916 41020 23660 41076
rect 23716 41020 23726 41076
rect 28466 41020 28476 41076
rect 28532 41020 29316 41076
rect 29698 41020 29708 41076
rect 29764 41020 29932 41076
rect 29988 41020 29998 41076
rect 30370 41020 30380 41076
rect 30436 41020 33852 41076
rect 33908 41020 33918 41076
rect 34748 41020 38332 41076
rect 38388 41020 38398 41076
rect 38612 41020 40124 41076
rect 40180 41020 40190 41076
rect 9212 40964 9268 41020
rect 29260 40964 29316 41020
rect 38612 40964 38668 41020
rect 49200 40992 49800 41104
rect 1922 40908 1932 40964
rect 1988 40908 7532 40964
rect 7588 40908 7598 40964
rect 7858 40908 7868 40964
rect 7924 40908 9268 40964
rect 13794 40908 13804 40964
rect 13860 40908 28812 40964
rect 28868 40908 28878 40964
rect 29260 40908 30268 40964
rect 30324 40908 31500 40964
rect 31556 40908 31566 40964
rect 32274 40908 32284 40964
rect 32340 40908 32396 40964
rect 32452 40908 32462 40964
rect 32610 40908 32620 40964
rect 32676 40908 32732 40964
rect 32788 40908 32798 40964
rect 33142 40908 33180 40964
rect 33236 40908 33246 40964
rect 33618 40908 33628 40964
rect 33684 40908 34972 40964
rect 35028 40908 35038 40964
rect 35522 40908 35532 40964
rect 35588 40908 35700 40964
rect 36390 40908 36428 40964
rect 36484 40908 36494 40964
rect 37398 40908 37436 40964
rect 37492 40908 37502 40964
rect 37874 40908 37884 40964
rect 37940 40908 38668 40964
rect 38994 40908 39004 40964
rect 39060 40908 39228 40964
rect 39284 40908 39294 40964
rect 35644 40852 35700 40908
rect 5058 40796 5068 40852
rect 5124 40796 8876 40852
rect 8932 40796 8942 40852
rect 9426 40796 9436 40852
rect 9492 40796 10444 40852
rect 10500 40796 10510 40852
rect 13458 40796 13468 40852
rect 13524 40796 16716 40852
rect 16772 40796 19628 40852
rect 19684 40796 19694 40852
rect 26450 40796 26460 40852
rect 26516 40796 35420 40852
rect 35476 40796 35486 40852
rect 35634 40796 35644 40852
rect 35700 40796 37100 40852
rect 37156 40796 37166 40852
rect 13468 40740 13524 40796
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 3938 40684 3948 40740
rect 4004 40684 6860 40740
rect 6916 40684 6926 40740
rect 7186 40684 7196 40740
rect 7252 40684 7420 40740
rect 7476 40684 7756 40740
rect 7812 40684 7822 40740
rect 7970 40684 7980 40740
rect 8036 40684 13524 40740
rect 16706 40684 16716 40740
rect 16772 40684 17612 40740
rect 17668 40684 17678 40740
rect 20972 40684 23436 40740
rect 23492 40684 23502 40740
rect 24546 40684 24556 40740
rect 24612 40684 29260 40740
rect 29316 40684 29326 40740
rect 29474 40684 29484 40740
rect 29540 40684 30380 40740
rect 30436 40684 33740 40740
rect 33796 40684 33806 40740
rect 34290 40684 34300 40740
rect 34356 40684 34860 40740
rect 34916 40684 34926 40740
rect 35186 40684 35196 40740
rect 35252 40684 37884 40740
rect 37940 40684 37950 40740
rect 20972 40628 21028 40684
rect 3490 40572 3500 40628
rect 3556 40572 9884 40628
rect 9940 40572 9950 40628
rect 13458 40572 13468 40628
rect 13524 40572 21028 40628
rect 21186 40572 21196 40628
rect 21252 40572 21420 40628
rect 21476 40572 21486 40628
rect 29362 40572 29372 40628
rect 29428 40572 29596 40628
rect 29652 40572 29662 40628
rect 31602 40572 31612 40628
rect 31668 40572 33404 40628
rect 33460 40572 33470 40628
rect 33618 40572 33628 40628
rect 33684 40572 38220 40628
rect 38276 40572 38286 40628
rect 3042 40460 3052 40516
rect 3108 40460 8428 40516
rect 8484 40460 13356 40516
rect 13412 40460 13422 40516
rect 13570 40460 13580 40516
rect 13636 40460 15932 40516
rect 15988 40460 15998 40516
rect 18060 40460 20188 40516
rect 20244 40460 20254 40516
rect 20402 40460 20412 40516
rect 20468 40460 22204 40516
rect 22260 40460 28028 40516
rect 28084 40460 28094 40516
rect 29474 40460 29484 40516
rect 29540 40460 30044 40516
rect 30100 40460 30110 40516
rect 30492 40460 31388 40516
rect 31444 40460 31454 40516
rect 31826 40460 31836 40516
rect 31892 40460 32284 40516
rect 32340 40460 32350 40516
rect 32498 40460 32508 40516
rect 32564 40460 32732 40516
rect 32788 40460 32798 40516
rect 32946 40460 32956 40516
rect 33012 40460 38668 40516
rect 38724 40460 38734 40516
rect 200 40320 800 40432
rect 18060 40404 18116 40460
rect 30492 40404 30548 40460
rect 2370 40348 2380 40404
rect 2436 40348 4060 40404
rect 4116 40348 4126 40404
rect 4386 40348 4396 40404
rect 4452 40348 9380 40404
rect 9622 40348 9660 40404
rect 9716 40348 9726 40404
rect 9874 40348 9884 40404
rect 9940 40348 9950 40404
rect 12002 40348 12012 40404
rect 12068 40348 14812 40404
rect 14868 40348 14878 40404
rect 15698 40348 15708 40404
rect 15764 40348 18060 40404
rect 18116 40348 18126 40404
rect 18274 40348 18284 40404
rect 18340 40348 18378 40404
rect 18498 40348 18508 40404
rect 18564 40348 20748 40404
rect 20804 40348 21532 40404
rect 21588 40348 21598 40404
rect 24406 40348 24444 40404
rect 24500 40348 24510 40404
rect 25106 40348 25116 40404
rect 25172 40348 30548 40404
rect 30902 40348 30940 40404
rect 30996 40348 31006 40404
rect 31164 40348 32620 40404
rect 32676 40348 32686 40404
rect 33058 40348 33068 40404
rect 33124 40348 33964 40404
rect 34020 40348 34030 40404
rect 34178 40348 34188 40404
rect 34244 40348 35644 40404
rect 35700 40348 35710 40404
rect 36194 40348 36204 40404
rect 36260 40348 36428 40404
rect 36484 40348 36494 40404
rect 38770 40348 38780 40404
rect 38836 40348 39116 40404
rect 39172 40348 39182 40404
rect 3602 40236 3612 40292
rect 3668 40236 6972 40292
rect 7028 40236 8876 40292
rect 8932 40236 8942 40292
rect 9324 40180 9380 40348
rect 9884 40292 9940 40348
rect 31164 40292 31220 40348
rect 9884 40236 11004 40292
rect 11060 40236 11070 40292
rect 13570 40236 13580 40292
rect 13636 40236 13916 40292
rect 13972 40236 13982 40292
rect 18946 40236 18956 40292
rect 19012 40236 20524 40292
rect 20580 40236 20590 40292
rect 22642 40236 22652 40292
rect 22708 40236 22988 40292
rect 23044 40236 23054 40292
rect 26450 40236 26460 40292
rect 26516 40236 29372 40292
rect 29428 40236 29438 40292
rect 29586 40236 29596 40292
rect 29652 40236 29708 40292
rect 29764 40236 29774 40292
rect 30258 40236 30268 40292
rect 30324 40236 31220 40292
rect 31836 40236 33740 40292
rect 33796 40236 33806 40292
rect 34402 40236 34412 40292
rect 34468 40236 37884 40292
rect 37940 40236 37950 40292
rect 31836 40180 31892 40236
rect 38612 40180 38668 40292
rect 38724 40236 38734 40292
rect 6066 40124 6076 40180
rect 6132 40124 6636 40180
rect 6692 40124 7756 40180
rect 7812 40124 7822 40180
rect 8614 40124 8652 40180
rect 8708 40124 8718 40180
rect 9324 40124 11340 40180
rect 11396 40124 11406 40180
rect 19170 40124 19180 40180
rect 19236 40124 20412 40180
rect 20468 40124 20478 40180
rect 25330 40124 25340 40180
rect 25396 40124 25788 40180
rect 25844 40124 27916 40180
rect 27972 40124 27982 40180
rect 29250 40124 29260 40180
rect 29316 40124 29820 40180
rect 29876 40124 31892 40180
rect 32050 40124 32060 40180
rect 32116 40124 32284 40180
rect 32340 40124 32350 40180
rect 32498 40124 32508 40180
rect 32564 40124 32732 40180
rect 32788 40124 38668 40180
rect 7830 40012 7868 40068
rect 7924 40012 7934 40068
rect 11778 40012 11788 40068
rect 11844 40012 22764 40068
rect 22820 40012 22830 40068
rect 26786 40012 26796 40068
rect 26852 40012 28700 40068
rect 28756 40012 31388 40068
rect 31444 40012 31500 40068
rect 31556 40012 31566 40068
rect 33058 40012 33068 40068
rect 33124 40012 34412 40068
rect 34468 40012 34478 40068
rect 34626 40012 34636 40068
rect 34692 40012 34860 40068
rect 34916 40012 34926 40068
rect 35532 40012 41468 40068
rect 41524 40012 41534 40068
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 5618 39900 5628 39956
rect 5684 39900 5694 39956
rect 6178 39900 6188 39956
rect 6244 39900 14644 39956
rect 15026 39900 15036 39956
rect 15092 39900 20300 39956
rect 20356 39900 21196 39956
rect 21252 39900 21262 39956
rect 21746 39900 21756 39956
rect 21812 39900 25228 39956
rect 25284 39900 25294 39956
rect 27234 39900 27244 39956
rect 27300 39900 28028 39956
rect 28084 39900 28094 39956
rect 29810 39900 29820 39956
rect 29876 39900 29932 39956
rect 29988 39900 29998 39956
rect 32498 39900 32508 39956
rect 32564 39900 33292 39956
rect 33348 39900 33358 39956
rect 33730 39900 33740 39956
rect 33796 39900 34412 39956
rect 34468 39900 34478 39956
rect 5628 39732 5684 39900
rect 14588 39844 14644 39900
rect 35532 39844 35588 40012
rect 35746 39900 35756 39956
rect 35812 39900 37100 39956
rect 37156 39900 37166 39956
rect 5842 39788 5852 39844
rect 5908 39788 9100 39844
rect 9156 39788 9166 39844
rect 10098 39788 10108 39844
rect 10164 39788 10556 39844
rect 10612 39788 10622 39844
rect 12338 39788 12348 39844
rect 12404 39788 12908 39844
rect 12964 39788 12974 39844
rect 14588 39788 16492 39844
rect 16548 39788 16558 39844
rect 19282 39788 19292 39844
rect 19348 39788 30044 39844
rect 30100 39788 30110 39844
rect 30258 39788 30268 39844
rect 30324 39788 30604 39844
rect 30660 39788 30670 39844
rect 30818 39788 30828 39844
rect 30884 39788 35084 39844
rect 35140 39788 35150 39844
rect 35298 39788 35308 39844
rect 35364 39788 35588 39844
rect 49200 39732 49800 39760
rect 2818 39676 2828 39732
rect 2884 39676 3612 39732
rect 3668 39676 3678 39732
rect 4498 39676 4508 39732
rect 4564 39676 5068 39732
rect 5124 39676 6860 39732
rect 6916 39676 6926 39732
rect 7410 39676 7420 39732
rect 7476 39676 18284 39732
rect 18340 39676 18350 39732
rect 20850 39676 20860 39732
rect 20916 39676 21644 39732
rect 21700 39676 21710 39732
rect 27122 39676 27132 39732
rect 27188 39676 30268 39732
rect 30324 39676 30334 39732
rect 30594 39676 30604 39732
rect 30660 39676 31164 39732
rect 31220 39676 31230 39732
rect 31938 39676 31948 39732
rect 32004 39676 32732 39732
rect 32788 39676 32798 39732
rect 33170 39676 33180 39732
rect 33236 39676 38668 39732
rect 48066 39676 48076 39732
rect 48132 39676 49800 39732
rect 33628 39620 33684 39676
rect 38612 39620 38668 39676
rect 49200 39648 49800 39676
rect 3266 39564 3276 39620
rect 3332 39564 7644 39620
rect 7700 39564 7710 39620
rect 9762 39564 9772 39620
rect 9828 39564 13916 39620
rect 13972 39564 13982 39620
rect 14466 39564 14476 39620
rect 14532 39564 15036 39620
rect 15092 39564 15102 39620
rect 17826 39564 17836 39620
rect 17892 39564 24556 39620
rect 24612 39564 24622 39620
rect 24770 39564 24780 39620
rect 24836 39564 26684 39620
rect 26740 39564 26750 39620
rect 28130 39564 28140 39620
rect 28196 39564 28476 39620
rect 28532 39564 30716 39620
rect 30772 39564 33292 39620
rect 33348 39564 33358 39620
rect 33590 39564 33628 39620
rect 33684 39564 33694 39620
rect 33842 39564 33852 39620
rect 33908 39564 38332 39620
rect 38388 39564 38398 39620
rect 38612 39564 38780 39620
rect 38836 39564 38846 39620
rect 6524 39452 10780 39508
rect 10836 39452 12460 39508
rect 12516 39452 12526 39508
rect 13542 39452 13580 39508
rect 13636 39452 13646 39508
rect 18694 39452 18732 39508
rect 18788 39452 18798 39508
rect 24434 39452 24444 39508
rect 24500 39452 24892 39508
rect 24948 39452 24958 39508
rect 27234 39452 27244 39508
rect 27300 39452 35084 39508
rect 35140 39452 35150 39508
rect 5404 39340 5852 39396
rect 5908 39340 5918 39396
rect 5404 39284 5460 39340
rect 4162 39228 4172 39284
rect 4228 39228 5404 39284
rect 5460 39228 5470 39284
rect 6524 39172 6580 39452
rect 6850 39340 6860 39396
rect 6916 39340 7420 39396
rect 7476 39340 7486 39396
rect 7634 39340 7644 39396
rect 7700 39340 8204 39396
rect 8260 39340 8270 39396
rect 8754 39340 8764 39396
rect 8820 39340 9100 39396
rect 9156 39340 9166 39396
rect 9398 39340 9436 39396
rect 9492 39340 9502 39396
rect 10210 39340 10220 39396
rect 10276 39340 10892 39396
rect 10948 39340 10958 39396
rect 13468 39340 20636 39396
rect 20692 39340 20702 39396
rect 21186 39340 21196 39396
rect 21252 39340 27468 39396
rect 27524 39340 27534 39396
rect 28690 39340 28700 39396
rect 28756 39340 28766 39396
rect 29250 39340 29260 39396
rect 29316 39340 29372 39396
rect 29428 39340 29438 39396
rect 29596 39340 30268 39396
rect 30324 39340 30334 39396
rect 30482 39340 30492 39396
rect 30548 39340 30558 39396
rect 31714 39340 31724 39396
rect 31780 39340 34748 39396
rect 34804 39340 34814 39396
rect 34972 39340 36092 39396
rect 36148 39340 36158 39396
rect 13468 39284 13524 39340
rect 20636 39284 20692 39340
rect 28700 39284 28756 39340
rect 29596 39284 29652 39340
rect 30492 39284 30548 39340
rect 34972 39284 35028 39340
rect 7792 39228 7868 39284
rect 7924 39228 13524 39284
rect 13794 39228 13804 39284
rect 13860 39228 15372 39284
rect 15428 39228 15438 39284
rect 20636 39228 27916 39284
rect 27972 39228 29652 39284
rect 29810 39228 29820 39284
rect 29876 39228 33292 39284
rect 33348 39228 33358 39284
rect 33478 39228 33516 39284
rect 33572 39228 33582 39284
rect 33730 39228 33740 39284
rect 33796 39228 34300 39284
rect 34356 39228 34366 39284
rect 34524 39228 35028 39284
rect 35186 39228 35196 39284
rect 35252 39228 35812 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 34524 39172 34580 39228
rect 2482 39116 2492 39172
rect 2548 39116 5852 39172
rect 5908 39116 6356 39172
rect 6514 39116 6524 39172
rect 6580 39116 6590 39172
rect 6748 39116 9772 39172
rect 9828 39116 9838 39172
rect 9986 39116 9996 39172
rect 10052 39116 18844 39172
rect 18900 39116 19180 39172
rect 19236 39116 19246 39172
rect 24546 39116 24556 39172
rect 24612 39116 31276 39172
rect 31332 39116 31836 39172
rect 31892 39116 31902 39172
rect 32386 39116 32396 39172
rect 32452 39116 32844 39172
rect 32900 39116 32910 39172
rect 33282 39116 33292 39172
rect 33348 39116 34580 39172
rect 34738 39116 34748 39172
rect 34804 39116 35420 39172
rect 35476 39116 35486 39172
rect 6300 39060 6356 39116
rect 6748 39060 6804 39116
rect 35756 39060 35812 39228
rect 35980 39116 36652 39172
rect 36708 39116 36718 39172
rect 35980 39060 36036 39116
rect 5058 39004 5068 39060
rect 5124 39004 6076 39060
rect 6132 39004 6142 39060
rect 6300 39004 6804 39060
rect 7746 39004 7756 39060
rect 7812 39004 9212 39060
rect 9268 39004 9772 39060
rect 9828 39004 9838 39060
rect 10518 39004 10556 39060
rect 10612 39004 10622 39060
rect 14018 39004 14028 39060
rect 14084 39004 27244 39060
rect 27300 39004 27310 39060
rect 27804 39004 32732 39060
rect 32788 39004 32798 39060
rect 33394 39004 33404 39060
rect 33460 39004 35532 39060
rect 35588 39004 35598 39060
rect 35756 39004 36036 39060
rect 36194 39004 36204 39060
rect 36260 39004 40908 39060
rect 40964 39004 40974 39060
rect 27804 38948 27860 39004
rect 6402 38892 6412 38948
rect 6468 38892 10108 38948
rect 10164 38892 10174 38948
rect 10322 38892 10332 38948
rect 10388 38892 12908 38948
rect 12964 38892 17164 38948
rect 17220 38892 17230 38948
rect 24658 38892 24668 38948
rect 24724 38892 25788 38948
rect 25844 38892 25854 38948
rect 27766 38892 27804 38948
rect 27860 38892 27870 38948
rect 28774 38892 28812 38948
rect 28868 38892 28878 38948
rect 29250 38892 29260 38948
rect 29316 38892 30156 38948
rect 30212 38892 30222 38948
rect 30370 38892 30380 38948
rect 30436 38892 30492 38948
rect 30548 38892 30558 38948
rect 31042 38892 31052 38948
rect 31108 38892 31164 38948
rect 31220 38892 31230 38948
rect 32162 38892 32172 38948
rect 32228 38892 32956 38948
rect 33012 38892 33022 38948
rect 34178 38892 34188 38948
rect 34244 38892 36316 38948
rect 36372 38892 37548 38948
rect 37604 38892 37614 38948
rect 4162 38780 4172 38836
rect 4228 38780 5740 38836
rect 5796 38780 8428 38836
rect 8484 38780 10220 38836
rect 10276 38780 13020 38836
rect 13076 38780 13086 38836
rect 13906 38780 13916 38836
rect 13972 38780 18844 38836
rect 18900 38780 18910 38836
rect 19618 38780 19628 38836
rect 19684 38780 25676 38836
rect 25732 38780 25742 38836
rect 27906 38780 27916 38836
rect 27972 38780 28476 38836
rect 28532 38780 28542 38836
rect 30034 38780 30044 38836
rect 30100 38780 30212 38836
rect 30370 38780 30380 38836
rect 30436 38780 32228 38836
rect 32386 38780 32396 38836
rect 32452 38780 32462 38836
rect 33058 38780 33068 38836
rect 33124 38780 33516 38836
rect 33572 38780 33582 38836
rect 33842 38780 33852 38836
rect 33908 38780 33964 38836
rect 34020 38780 35084 38836
rect 35140 38780 35150 38836
rect 35298 38780 35308 38836
rect 35364 38780 38668 38836
rect 38724 38780 40012 38836
rect 40068 38780 40078 38836
rect 30156 38724 30212 38780
rect 5506 38668 5516 38724
rect 5572 38668 6524 38724
rect 6580 38668 6590 38724
rect 7298 38668 7308 38724
rect 7364 38668 7420 38724
rect 7476 38668 7486 38724
rect 7746 38668 7756 38724
rect 7812 38668 7980 38724
rect 8036 38668 10332 38724
rect 10388 38668 10398 38724
rect 10546 38668 10556 38724
rect 10612 38668 12684 38724
rect 12740 38668 12750 38724
rect 13234 38668 13244 38724
rect 13300 38668 13356 38724
rect 13412 38668 13422 38724
rect 13916 38668 19852 38724
rect 19908 38668 19918 38724
rect 21858 38668 21868 38724
rect 21924 38668 24276 38724
rect 24434 38668 24444 38724
rect 24500 38668 24556 38724
rect 24612 38668 24622 38724
rect 24780 38668 24892 38724
rect 24948 38668 25396 38724
rect 26338 38668 26348 38724
rect 26404 38668 26908 38724
rect 26964 38668 26974 38724
rect 28018 38668 28028 38724
rect 28084 38668 30100 38724
rect 30156 38668 31948 38724
rect 32004 38668 32014 38724
rect 13916 38612 13972 38668
rect 24220 38612 24276 38668
rect 24780 38612 24836 38668
rect 3332 38556 12516 38612
rect 12674 38556 12684 38612
rect 12740 38556 13972 38612
rect 15362 38556 15372 38612
rect 15428 38556 16156 38612
rect 16212 38556 19516 38612
rect 19572 38556 19582 38612
rect 21634 38556 21644 38612
rect 21700 38556 21980 38612
rect 22036 38556 22316 38612
rect 22372 38556 22382 38612
rect 24220 38556 24836 38612
rect 25340 38612 25396 38668
rect 30044 38612 30100 38668
rect 32172 38612 32228 38780
rect 32396 38724 32452 38780
rect 32396 38668 32508 38724
rect 32564 38668 36092 38724
rect 36148 38668 36158 38724
rect 25340 38556 28700 38612
rect 28756 38556 28766 38612
rect 30034 38556 30044 38612
rect 30100 38556 30110 38612
rect 30258 38556 30268 38612
rect 30324 38556 32004 38612
rect 32172 38556 34076 38612
rect 34132 38556 34300 38612
rect 34356 38556 34366 38612
rect 34524 38556 35980 38612
rect 36036 38556 36046 38612
rect 36530 38556 36540 38612
rect 36596 38556 39452 38612
rect 39508 38556 39518 38612
rect 200 38388 800 38416
rect 200 38332 1820 38388
rect 1876 38332 1886 38388
rect 200 38304 800 38332
rect 3332 38276 3388 38556
rect 12460 38500 12516 38556
rect 31948 38500 32004 38556
rect 34524 38500 34580 38556
rect 5628 38444 11116 38500
rect 11172 38444 11452 38500
rect 11508 38444 11518 38500
rect 11666 38444 11676 38500
rect 11732 38444 12236 38500
rect 12292 38444 12302 38500
rect 12460 38444 12572 38500
rect 12628 38444 14364 38500
rect 14420 38444 14430 38500
rect 25890 38444 25900 38500
rect 25956 38444 28700 38500
rect 28756 38444 28766 38500
rect 30370 38444 30380 38500
rect 30436 38444 31052 38500
rect 31108 38444 31118 38500
rect 31266 38444 31276 38500
rect 31332 38444 31724 38500
rect 31780 38444 31790 38500
rect 31938 38444 31948 38500
rect 32004 38444 34580 38500
rect 35830 38444 35868 38500
rect 35924 38444 35934 38500
rect 36092 38444 37324 38500
rect 37380 38444 37390 38500
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 5628 38276 5684 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 5842 38332 5852 38388
rect 5908 38332 11004 38388
rect 11060 38332 11340 38388
rect 11396 38332 11406 38388
rect 12002 38332 12012 38388
rect 12068 38332 15148 38388
rect 17042 38332 17052 38388
rect 17108 38332 27580 38388
rect 27636 38332 27646 38388
rect 30258 38332 30268 38388
rect 30324 38332 31612 38388
rect 31668 38332 31678 38388
rect 31826 38332 31836 38388
rect 31892 38332 34524 38388
rect 34580 38332 34590 38388
rect 15092 38276 15148 38332
rect 36092 38276 36148 38444
rect 2930 38220 2940 38276
rect 2996 38220 3388 38276
rect 4610 38220 4620 38276
rect 4676 38220 5684 38276
rect 7410 38220 7420 38276
rect 7476 38220 11060 38276
rect 11218 38220 11228 38276
rect 11284 38220 13692 38276
rect 13748 38220 13758 38276
rect 15092 38220 16156 38276
rect 16212 38220 16222 38276
rect 18498 38220 18508 38276
rect 18564 38220 29708 38276
rect 29764 38220 29774 38276
rect 30146 38220 30156 38276
rect 30212 38220 30828 38276
rect 30884 38220 30894 38276
rect 31164 38220 31276 38276
rect 31332 38220 31342 38276
rect 31490 38220 31500 38276
rect 31556 38220 36148 38276
rect 11004 38164 11060 38220
rect 31164 38164 31220 38220
rect 4050 38108 4060 38164
rect 4116 38108 4956 38164
rect 5012 38108 8540 38164
rect 8596 38108 9996 38164
rect 10052 38108 10062 38164
rect 10658 38108 10668 38164
rect 10724 38108 10780 38164
rect 10836 38108 10846 38164
rect 11004 38108 13468 38164
rect 13524 38108 13534 38164
rect 14018 38108 14028 38164
rect 14084 38108 16492 38164
rect 16548 38108 16558 38164
rect 17378 38108 17388 38164
rect 17444 38108 17836 38164
rect 17892 38108 17902 38164
rect 18050 38108 18060 38164
rect 18116 38108 20860 38164
rect 20916 38108 22428 38164
rect 22484 38108 22494 38164
rect 26226 38108 26236 38164
rect 26292 38108 29148 38164
rect 29204 38108 29214 38164
rect 29474 38108 29484 38164
rect 29540 38108 31220 38164
rect 31276 38108 31724 38164
rect 31780 38108 31790 38164
rect 34290 38108 34300 38164
rect 34356 38108 34860 38164
rect 34916 38108 36540 38164
rect 36596 38108 36606 38164
rect 31276 38052 31332 38108
rect 6738 37996 6748 38052
rect 6804 37996 7588 38052
rect 7746 37996 7756 38052
rect 7812 37996 12404 38052
rect 12562 37996 12572 38052
rect 12628 37996 18284 38052
rect 18340 37996 18350 38052
rect 19058 37996 19068 38052
rect 19124 37996 19628 38052
rect 19684 37996 19694 38052
rect 20738 37996 20748 38052
rect 20804 37996 21644 38052
rect 21700 37996 21710 38052
rect 21868 37996 23324 38052
rect 23380 37996 23390 38052
rect 24098 37996 24108 38052
rect 24164 37996 28700 38052
rect 28756 37996 28766 38052
rect 28914 37996 28924 38052
rect 28980 37996 29036 38052
rect 29092 37996 31332 38052
rect 31490 37996 31500 38052
rect 31556 37996 32620 38052
rect 32676 37996 34636 38052
rect 34692 37996 34702 38052
rect 35746 37996 35756 38052
rect 35812 37996 35868 38052
rect 35924 37996 36764 38052
rect 36820 37996 36830 38052
rect 38612 37996 39564 38052
rect 39620 37996 39630 38052
rect 7532 37940 7588 37996
rect 12348 37940 12404 37996
rect 21868 37940 21924 37996
rect 5058 37884 5068 37940
rect 5124 37884 7308 37940
rect 7364 37884 7374 37940
rect 7522 37884 7532 37940
rect 7588 37884 8092 37940
rect 8148 37884 8428 37940
rect 8484 37884 9324 37940
rect 9380 37884 9390 37940
rect 10294 37884 10332 37940
rect 10388 37884 10398 37940
rect 10546 37884 10556 37940
rect 10612 37884 11116 37940
rect 11172 37884 11182 37940
rect 11330 37884 11340 37940
rect 11396 37884 12292 37940
rect 12348 37884 13692 37940
rect 13748 37884 14140 37940
rect 14196 37884 14206 37940
rect 18050 37884 18060 37940
rect 18116 37884 21868 37940
rect 21924 37884 21934 37940
rect 22418 37884 22428 37940
rect 22484 37884 25004 37940
rect 25060 37884 25070 37940
rect 29586 37884 29596 37940
rect 29652 37884 33964 37940
rect 34020 37884 34030 37940
rect 34822 37884 34860 37940
rect 34916 37884 34926 37940
rect 12236 37828 12292 37884
rect 7186 37772 7196 37828
rect 7252 37772 11900 37828
rect 11956 37772 11966 37828
rect 12236 37772 13244 37828
rect 13300 37772 13310 37828
rect 13458 37772 13468 37828
rect 13524 37772 15036 37828
rect 15092 37772 15102 37828
rect 18386 37772 18396 37828
rect 18452 37772 22092 37828
rect 22148 37772 22158 37828
rect 23426 37772 23436 37828
rect 23492 37772 25900 37828
rect 25956 37772 25966 37828
rect 27122 37772 27132 37828
rect 27188 37772 27468 37828
rect 27524 37772 27534 37828
rect 28662 37772 28700 37828
rect 28756 37772 28766 37828
rect 28914 37772 28924 37828
rect 28980 37772 29484 37828
rect 29540 37772 29550 37828
rect 29698 37772 29708 37828
rect 29764 37772 30044 37828
rect 30100 37772 30110 37828
rect 30258 37772 30268 37828
rect 30324 37772 30828 37828
rect 30884 37772 30894 37828
rect 31266 37772 31276 37828
rect 31332 37772 33180 37828
rect 33236 37772 35308 37828
rect 35364 37772 35374 37828
rect 35746 37772 35756 37828
rect 35812 37772 37100 37828
rect 37156 37772 37166 37828
rect 38612 37716 38668 37996
rect 49200 37716 49800 37744
rect 9986 37660 9996 37716
rect 10052 37660 18732 37716
rect 18788 37660 18956 37716
rect 19012 37660 19022 37716
rect 21970 37660 21980 37716
rect 22036 37660 22764 37716
rect 22820 37660 22830 37716
rect 28588 37660 33516 37716
rect 33572 37660 33740 37716
rect 33796 37660 33806 37716
rect 33954 37660 33964 37716
rect 34020 37660 38668 37716
rect 48066 37660 48076 37716
rect 48132 37660 49800 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 28588 37604 28644 37660
rect 49200 37632 49800 37660
rect 8642 37548 8652 37604
rect 8708 37548 12012 37604
rect 12068 37548 12078 37604
rect 12226 37548 12236 37604
rect 12292 37548 13804 37604
rect 13860 37548 14812 37604
rect 14868 37548 14878 37604
rect 22194 37548 22204 37604
rect 22260 37548 23884 37604
rect 23940 37548 25116 37604
rect 25172 37548 25182 37604
rect 25330 37548 25340 37604
rect 25396 37548 28588 37604
rect 28644 37548 28654 37604
rect 29026 37548 29036 37604
rect 29092 37548 29484 37604
rect 29540 37548 29708 37604
rect 29764 37548 29774 37604
rect 29922 37548 29932 37604
rect 29988 37548 36428 37604
rect 36484 37548 36494 37604
rect 5954 37436 5964 37492
rect 6020 37436 7868 37492
rect 7924 37436 7934 37492
rect 8764 37436 9884 37492
rect 9940 37436 9950 37492
rect 10210 37436 10220 37492
rect 10276 37436 11564 37492
rect 11620 37436 15148 37492
rect 19506 37436 19516 37492
rect 19572 37436 29596 37492
rect 29652 37436 29662 37492
rect 29820 37436 31500 37492
rect 31556 37436 34076 37492
rect 34132 37436 34142 37492
rect 34626 37436 34636 37492
rect 34692 37436 34860 37492
rect 34916 37436 34926 37492
rect 8764 37380 8820 37436
rect 15092 37380 15148 37436
rect 29820 37380 29876 37436
rect 2706 37324 2716 37380
rect 2772 37324 8764 37380
rect 8820 37324 8830 37380
rect 8950 37324 8988 37380
rect 9044 37324 9054 37380
rect 9986 37324 9996 37380
rect 10052 37324 10556 37380
rect 10612 37324 10622 37380
rect 10780 37324 12236 37380
rect 12292 37324 12302 37380
rect 13234 37324 13244 37380
rect 13300 37324 14028 37380
rect 14084 37324 14094 37380
rect 15092 37324 18956 37380
rect 19012 37324 19022 37380
rect 22530 37324 22540 37380
rect 22596 37324 25900 37380
rect 25956 37324 25966 37380
rect 27794 37324 27804 37380
rect 27860 37324 28588 37380
rect 28644 37324 28654 37380
rect 28802 37324 28812 37380
rect 28868 37324 29260 37380
rect 29316 37324 29876 37380
rect 30370 37324 30380 37380
rect 30436 37324 30492 37380
rect 30548 37324 33964 37380
rect 34020 37324 34030 37380
rect 34514 37324 34524 37380
rect 34580 37324 34748 37380
rect 34804 37324 34814 37380
rect 10780 37268 10836 37324
rect 14028 37268 14084 37324
rect 6850 37212 6860 37268
rect 6916 37212 10836 37268
rect 10994 37212 11004 37268
rect 11060 37212 12348 37268
rect 12404 37212 12414 37268
rect 14028 37212 15260 37268
rect 15316 37212 15326 37268
rect 16370 37212 16380 37268
rect 16436 37212 18396 37268
rect 18452 37212 20188 37268
rect 20244 37212 20254 37268
rect 21858 37212 21868 37268
rect 21924 37212 27020 37268
rect 27076 37212 28028 37268
rect 28084 37212 28094 37268
rect 28354 37212 28364 37268
rect 28420 37212 29708 37268
rect 29764 37212 29774 37268
rect 30034 37212 30044 37268
rect 30100 37212 33516 37268
rect 33572 37212 36876 37268
rect 36932 37212 36942 37268
rect 7186 37100 7196 37156
rect 7252 37100 7980 37156
rect 8036 37100 8046 37156
rect 8194 37100 8204 37156
rect 8260 37100 13468 37156
rect 13524 37100 21756 37156
rect 21812 37100 21822 37156
rect 22306 37100 22316 37156
rect 22372 37100 24444 37156
rect 24500 37100 25228 37156
rect 25284 37100 25294 37156
rect 26002 37100 26012 37156
rect 26068 37100 26236 37156
rect 26292 37100 26302 37156
rect 26852 37100 30940 37156
rect 30996 37100 31006 37156
rect 31602 37100 31612 37156
rect 31668 37100 32172 37156
rect 32228 37100 32238 37156
rect 32732 37100 33684 37156
rect 34402 37100 34412 37156
rect 34468 37100 36540 37156
rect 36596 37100 36606 37156
rect 200 37044 800 37072
rect 26852 37044 26908 37100
rect 32732 37044 32788 37100
rect 33628 37044 33684 37100
rect 200 36988 1820 37044
rect 1876 36988 1886 37044
rect 9314 36988 9324 37044
rect 9380 36988 9660 37044
rect 9716 36988 9726 37044
rect 9874 36988 9884 37044
rect 9940 36988 10276 37044
rect 10518 36988 10556 37044
rect 10612 36988 10622 37044
rect 10770 36988 10780 37044
rect 10836 36988 11788 37044
rect 11844 36988 16380 37044
rect 16436 36988 16446 37044
rect 16594 36988 16604 37044
rect 16660 36988 18060 37044
rect 18116 36988 18126 37044
rect 18386 36988 18396 37044
rect 18452 36988 22428 37044
rect 22484 36988 22494 37044
rect 23062 36988 23100 37044
rect 23156 36988 23166 37044
rect 24658 36988 24668 37044
rect 24724 36988 25340 37044
rect 25396 36988 25406 37044
rect 26114 36988 26124 37044
rect 26180 36988 26908 37044
rect 29810 36988 29820 37044
rect 29876 36988 30380 37044
rect 30436 36988 30446 37044
rect 30594 36988 30604 37044
rect 30660 36988 32788 37044
rect 32946 36988 32956 37044
rect 33012 36988 33404 37044
rect 33460 36988 33470 37044
rect 33628 36988 36204 37044
rect 36260 36988 36270 37044
rect 200 36960 800 36988
rect 10220 36932 10276 36988
rect 4834 36876 4844 36932
rect 4900 36876 9660 36932
rect 9716 36876 9726 36932
rect 10220 36876 12012 36932
rect 12068 36876 12078 36932
rect 14242 36876 14252 36932
rect 14308 36876 21868 36932
rect 21924 36876 21934 36932
rect 24210 36876 24220 36932
rect 24276 36876 27356 36932
rect 27412 36876 27422 36932
rect 28578 36876 28588 36932
rect 28644 36876 31724 36932
rect 31780 36876 31790 36932
rect 32582 36876 32620 36932
rect 32676 36876 32686 36932
rect 33842 36876 33852 36932
rect 33908 36876 34300 36932
rect 34356 36876 34366 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 5618 36764 5628 36820
rect 5684 36764 10108 36820
rect 10164 36764 10174 36820
rect 12012 36708 12068 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 12562 36764 12572 36820
rect 12628 36764 13356 36820
rect 13412 36764 17388 36820
rect 17444 36764 17454 36820
rect 17602 36764 17612 36820
rect 17668 36764 21980 36820
rect 22036 36764 22046 36820
rect 27682 36764 27692 36820
rect 27748 36764 28476 36820
rect 28532 36764 32732 36820
rect 32788 36764 32798 36820
rect 4834 36652 4844 36708
rect 4900 36652 11004 36708
rect 11060 36652 11070 36708
rect 12012 36652 12572 36708
rect 12628 36652 15372 36708
rect 15428 36652 15438 36708
rect 17276 36652 19292 36708
rect 19348 36652 20748 36708
rect 20804 36652 20814 36708
rect 24546 36652 24556 36708
rect 24612 36652 25228 36708
rect 25284 36652 25294 36708
rect 26002 36652 26012 36708
rect 26068 36652 30380 36708
rect 30436 36652 30446 36708
rect 30706 36652 30716 36708
rect 30772 36652 31612 36708
rect 31668 36652 31678 36708
rect 32274 36652 32284 36708
rect 32340 36652 38780 36708
rect 38836 36652 38846 36708
rect 17276 36596 17332 36652
rect 6290 36540 6300 36596
rect 6356 36540 6412 36596
rect 6468 36540 6478 36596
rect 8082 36540 8092 36596
rect 8148 36540 8428 36596
rect 8484 36540 8494 36596
rect 8866 36540 8876 36596
rect 8932 36540 13804 36596
rect 13860 36540 13870 36596
rect 14578 36540 14588 36596
rect 14644 36540 16828 36596
rect 16884 36540 17276 36596
rect 17332 36540 17342 36596
rect 17826 36540 17836 36596
rect 17892 36540 17948 36596
rect 18004 36540 18014 36596
rect 21634 36540 21644 36596
rect 21700 36540 21756 36596
rect 21812 36540 21822 36596
rect 23734 36540 23772 36596
rect 23828 36540 23838 36596
rect 26338 36540 26348 36596
rect 26404 36540 29932 36596
rect 29988 36540 29998 36596
rect 30146 36540 30156 36596
rect 30212 36540 30828 36596
rect 30884 36540 30894 36596
rect 31612 36484 31668 36652
rect 32162 36540 32172 36596
rect 32228 36540 39340 36596
rect 39396 36540 39406 36596
rect 6402 36428 6412 36484
rect 6468 36428 12572 36484
rect 12628 36428 12638 36484
rect 13990 36428 14028 36484
rect 14084 36428 14094 36484
rect 17724 36428 19516 36484
rect 19572 36428 20076 36484
rect 20132 36428 20142 36484
rect 20514 36428 20524 36484
rect 20580 36428 25340 36484
rect 25396 36428 25406 36484
rect 27122 36428 27132 36484
rect 27188 36428 30380 36484
rect 30436 36428 30446 36484
rect 31612 36428 35868 36484
rect 35924 36428 35934 36484
rect 17724 36372 17780 36428
rect 25340 36372 25396 36428
rect 9314 36316 9324 36372
rect 9380 36316 9772 36372
rect 9828 36316 9838 36372
rect 11218 36316 11228 36372
rect 11284 36316 17724 36372
rect 17780 36316 17790 36372
rect 17938 36316 17948 36372
rect 18004 36316 22988 36372
rect 23044 36316 23054 36372
rect 25340 36316 26012 36372
rect 26068 36316 26078 36372
rect 26758 36316 26796 36372
rect 26852 36316 26862 36372
rect 27234 36316 27244 36372
rect 27300 36316 31724 36372
rect 31780 36316 31790 36372
rect 31938 36316 31948 36372
rect 32004 36316 33516 36372
rect 33572 36316 33582 36372
rect 6710 36204 6748 36260
rect 6804 36204 8204 36260
rect 8260 36204 8270 36260
rect 8978 36204 8988 36260
rect 9044 36204 11676 36260
rect 11732 36204 11742 36260
rect 12002 36204 12012 36260
rect 12068 36204 12124 36260
rect 12180 36204 12190 36260
rect 12338 36204 12348 36260
rect 12404 36204 12908 36260
rect 12964 36204 13244 36260
rect 13300 36204 13310 36260
rect 13794 36204 13804 36260
rect 13860 36204 17724 36260
rect 17780 36204 17790 36260
rect 18946 36204 18956 36260
rect 19012 36204 28364 36260
rect 28420 36204 28430 36260
rect 28774 36204 28812 36260
rect 28868 36204 28878 36260
rect 29250 36204 29260 36260
rect 29316 36204 30044 36260
rect 30100 36204 30110 36260
rect 30706 36204 30716 36260
rect 30772 36204 31612 36260
rect 31668 36204 31678 36260
rect 31826 36204 31836 36260
rect 31892 36204 32844 36260
rect 32900 36204 32910 36260
rect 2594 36092 2604 36148
rect 2660 36092 8652 36148
rect 8708 36092 11788 36148
rect 11844 36092 12572 36148
rect 12628 36092 12638 36148
rect 13010 36092 13020 36148
rect 13076 36092 13692 36148
rect 13748 36092 13758 36148
rect 15026 36092 15036 36148
rect 15092 36092 18172 36148
rect 18228 36092 18238 36148
rect 25824 36092 25900 36148
rect 25956 36092 30604 36148
rect 30660 36092 30670 36148
rect 31266 36092 31276 36148
rect 31332 36092 32172 36148
rect 32228 36092 32238 36148
rect 32722 36092 32732 36148
rect 32788 36092 32956 36148
rect 33012 36092 35644 36148
rect 35700 36092 35710 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 5170 35980 5180 36036
rect 5236 35980 9996 36036
rect 10052 35980 10062 36036
rect 10368 35980 10444 36036
rect 10500 35980 12124 36036
rect 12180 35980 12190 36036
rect 12898 35980 12908 36036
rect 12964 35980 13132 36036
rect 13188 35980 18508 36036
rect 18564 35980 18574 36036
rect 27458 35980 27468 36036
rect 27524 35980 28028 36036
rect 28084 35980 28094 36036
rect 28242 35980 28252 36036
rect 28308 35980 31388 36036
rect 31444 35980 33068 36036
rect 33124 35980 33134 36036
rect 10770 35868 10780 35924
rect 10836 35868 11788 35924
rect 11844 35868 11854 35924
rect 14466 35868 14476 35924
rect 14532 35868 15708 35924
rect 15764 35868 15774 35924
rect 16594 35868 16604 35924
rect 16660 35868 27020 35924
rect 27076 35868 27086 35924
rect 27654 35868 27692 35924
rect 27748 35868 28476 35924
rect 28532 35868 28980 35924
rect 29110 35868 29148 35924
rect 29204 35868 29214 35924
rect 29372 35868 31276 35924
rect 31332 35868 31342 35924
rect 31602 35868 31612 35924
rect 31668 35868 31948 35924
rect 32004 35868 32014 35924
rect 28924 35812 28980 35868
rect 29372 35812 29428 35868
rect 9762 35756 9772 35812
rect 9828 35756 12460 35812
rect 12516 35756 12526 35812
rect 15026 35756 15036 35812
rect 15092 35756 17724 35812
rect 17780 35756 17790 35812
rect 17938 35756 17948 35812
rect 18004 35756 18172 35812
rect 18228 35756 18238 35812
rect 18498 35756 18508 35812
rect 18564 35756 20076 35812
rect 20132 35756 20142 35812
rect 23090 35756 23100 35812
rect 23156 35756 24220 35812
rect 24276 35756 24780 35812
rect 24836 35756 24846 35812
rect 28550 35756 28588 35812
rect 28644 35756 28654 35812
rect 28924 35756 29428 35812
rect 29586 35756 29596 35812
rect 29652 35756 32396 35812
rect 32452 35756 32462 35812
rect 49200 35700 49800 35728
rect 8642 35644 8652 35700
rect 8708 35644 11116 35700
rect 11172 35644 11182 35700
rect 13458 35644 13468 35700
rect 13524 35644 15036 35700
rect 15092 35644 15102 35700
rect 15586 35644 15596 35700
rect 15652 35644 16044 35700
rect 16100 35644 16110 35700
rect 16930 35644 16940 35700
rect 16996 35644 21084 35700
rect 21140 35644 21150 35700
rect 25218 35644 25228 35700
rect 25284 35644 25676 35700
rect 25732 35644 25742 35700
rect 26124 35644 31500 35700
rect 31556 35644 31566 35700
rect 31714 35644 31724 35700
rect 31780 35644 33628 35700
rect 33684 35644 33694 35700
rect 48066 35644 48076 35700
rect 48132 35644 49800 35700
rect 7270 35532 7308 35588
rect 7364 35532 7374 35588
rect 7746 35532 7756 35588
rect 7812 35532 9100 35588
rect 9156 35532 9166 35588
rect 10210 35532 10220 35588
rect 10276 35532 10286 35588
rect 11666 35532 11676 35588
rect 11732 35532 18340 35588
rect 18498 35532 18508 35588
rect 18564 35532 24332 35588
rect 24388 35532 24398 35588
rect 24882 35532 24892 35588
rect 24948 35532 25676 35588
rect 25732 35532 25742 35588
rect 10220 35476 10276 35532
rect 18284 35476 18340 35532
rect 26124 35476 26180 35644
rect 49200 35616 49800 35644
rect 27318 35532 27356 35588
rect 27412 35532 27422 35588
rect 27570 35532 27580 35588
rect 27636 35532 27692 35588
rect 27748 35532 29652 35588
rect 29810 35532 29820 35588
rect 29876 35532 39004 35588
rect 39060 35532 39070 35588
rect 29596 35476 29652 35532
rect 10220 35420 12012 35476
rect 12068 35420 14364 35476
rect 14420 35420 14430 35476
rect 15092 35420 16604 35476
rect 16660 35420 16670 35476
rect 17490 35420 17500 35476
rect 17556 35420 17948 35476
rect 18004 35420 18014 35476
rect 18284 35420 18396 35476
rect 18452 35420 18462 35476
rect 20178 35420 20188 35476
rect 20244 35420 25396 35476
rect 26086 35420 26124 35476
rect 26180 35420 26190 35476
rect 26348 35420 27132 35476
rect 27188 35420 27198 35476
rect 27356 35420 29540 35476
rect 29596 35420 29708 35476
rect 29764 35420 32732 35476
rect 32788 35420 32798 35476
rect 15092 35364 15148 35420
rect 25340 35364 25396 35420
rect 26348 35364 26404 35420
rect 27356 35364 27412 35420
rect 29484 35364 29540 35420
rect 5618 35308 5628 35364
rect 5684 35308 6524 35364
rect 6580 35308 6590 35364
rect 11788 35308 15148 35364
rect 15586 35308 15596 35364
rect 15652 35308 23828 35364
rect 23986 35308 23996 35364
rect 24052 35308 25116 35364
rect 25172 35308 25182 35364
rect 25340 35308 26404 35364
rect 26562 35308 26572 35364
rect 26628 35308 27412 35364
rect 27570 35308 27580 35364
rect 27636 35308 29316 35364
rect 29474 35308 29484 35364
rect 29540 35308 29596 35364
rect 29652 35308 29662 35364
rect 29820 35308 30156 35364
rect 30212 35308 30222 35364
rect 30790 35308 30828 35364
rect 30884 35308 30894 35364
rect 32162 35308 32172 35364
rect 32228 35308 33068 35364
rect 33124 35308 33134 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 11788 35252 11844 35308
rect 23772 35252 23828 35308
rect 29260 35252 29316 35308
rect 29820 35252 29876 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 9538 35196 9548 35252
rect 9604 35196 11844 35252
rect 13682 35196 13692 35252
rect 13748 35196 13804 35252
rect 13860 35196 13870 35252
rect 14886 35196 14924 35252
rect 14980 35196 14990 35252
rect 17378 35196 17388 35252
rect 17444 35196 23548 35252
rect 23604 35196 23614 35252
rect 23772 35196 25284 35252
rect 25442 35196 25452 35252
rect 25508 35196 27412 35252
rect 27682 35196 27692 35252
rect 27748 35196 27916 35252
rect 27972 35196 27982 35252
rect 28242 35196 28252 35252
rect 28308 35196 28476 35252
rect 28532 35196 28542 35252
rect 29260 35196 29876 35252
rect 30930 35196 30940 35252
rect 30996 35196 31164 35252
rect 31220 35196 31230 35252
rect 32722 35196 32732 35252
rect 32788 35196 33964 35252
rect 34020 35196 34030 35252
rect 10332 35140 10388 35196
rect 25228 35140 25284 35196
rect 27356 35140 27412 35196
rect 10322 35084 10332 35140
rect 10388 35084 10398 35140
rect 11554 35084 11564 35140
rect 11620 35084 15820 35140
rect 15876 35084 16492 35140
rect 16548 35084 16558 35140
rect 21746 35084 21756 35140
rect 21812 35084 21980 35140
rect 22036 35084 22046 35140
rect 25228 35084 27020 35140
rect 27076 35084 27086 35140
rect 27346 35084 27356 35140
rect 27412 35084 29932 35140
rect 29988 35084 29998 35140
rect 31266 35084 31276 35140
rect 31332 35084 38556 35140
rect 38612 35084 38622 35140
rect 200 35028 800 35056
rect 200 34972 1820 35028
rect 1876 34972 1886 35028
rect 7074 34972 7084 35028
rect 7140 34972 8204 35028
rect 8260 34972 8876 35028
rect 8932 34972 8942 35028
rect 15036 34972 17388 35028
rect 17444 34972 17454 35028
rect 18274 34972 18284 35028
rect 18340 34972 21644 35028
rect 21700 34972 21710 35028
rect 22418 34972 22428 35028
rect 22484 34972 23884 35028
rect 23940 34972 23950 35028
rect 24210 34972 24220 35028
rect 24276 34972 30940 35028
rect 30996 34972 31006 35028
rect 200 34944 800 34972
rect 15036 34916 15092 34972
rect 11218 34860 11228 34916
rect 11284 34860 12684 34916
rect 12740 34860 15092 34916
rect 21634 34860 21644 34916
rect 21700 34860 26908 34916
rect 28578 34860 28588 34916
rect 28644 34860 30492 34916
rect 30548 34860 32284 34916
rect 32340 34860 32350 34916
rect 26852 34804 26908 34860
rect 10994 34748 11004 34804
rect 11060 34748 13804 34804
rect 13860 34748 13870 34804
rect 14662 34748 14700 34804
rect 14756 34748 14766 34804
rect 16258 34748 16268 34804
rect 16324 34748 16380 34804
rect 16436 34748 16446 34804
rect 18498 34748 18508 34804
rect 18564 34748 20076 34804
rect 20132 34748 20142 34804
rect 23538 34748 23548 34804
rect 23604 34748 23772 34804
rect 23828 34748 23838 34804
rect 25106 34748 25116 34804
rect 25172 34748 25788 34804
rect 25844 34748 25854 34804
rect 26852 34748 27020 34804
rect 27076 34748 32396 34804
rect 32452 34748 32462 34804
rect 9874 34636 9884 34692
rect 9940 34636 10668 34692
rect 10724 34636 10734 34692
rect 11218 34636 11228 34692
rect 11284 34636 12572 34692
rect 12628 34636 12638 34692
rect 15922 34636 15932 34692
rect 15988 34636 25004 34692
rect 25060 34636 25070 34692
rect 25218 34636 25228 34692
rect 25284 34636 27916 34692
rect 27972 34636 27982 34692
rect 32162 34636 32172 34692
rect 32228 34636 34972 34692
rect 35028 34636 35038 34692
rect 5282 34524 5292 34580
rect 5348 34524 11564 34580
rect 11620 34524 11630 34580
rect 12114 34524 12124 34580
rect 12180 34524 15820 34580
rect 15876 34524 16156 34580
rect 16212 34524 16222 34580
rect 16370 34524 16380 34580
rect 16436 34524 16492 34580
rect 16548 34524 16558 34580
rect 17378 34524 17388 34580
rect 17444 34524 18564 34580
rect 23874 34524 23884 34580
rect 23940 34524 25900 34580
rect 25956 34524 25966 34580
rect 26852 34524 30380 34580
rect 30436 34524 35868 34580
rect 35924 34524 35934 34580
rect 11564 34468 11620 34524
rect 9426 34412 9436 34468
rect 9492 34412 11004 34468
rect 11060 34412 11070 34468
rect 11564 34412 13468 34468
rect 13524 34412 13534 34468
rect 13682 34412 13692 34468
rect 13748 34412 16716 34468
rect 16772 34412 18284 34468
rect 18340 34412 18350 34468
rect 18508 34356 18564 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 26852 34468 26908 34524
rect 26002 34412 26012 34468
rect 26068 34412 26908 34468
rect 27122 34412 27132 34468
rect 27188 34412 27580 34468
rect 27636 34412 28476 34468
rect 28532 34412 35532 34468
rect 35588 34412 35598 34468
rect 49200 34356 49800 34384
rect 8754 34300 8764 34356
rect 8820 34300 12460 34356
rect 12516 34300 12526 34356
rect 14242 34300 14252 34356
rect 14308 34300 14924 34356
rect 14980 34300 14990 34356
rect 15082 34300 15092 34356
rect 15148 34300 18060 34356
rect 18116 34300 18126 34356
rect 18508 34300 20860 34356
rect 20916 34300 20926 34356
rect 22540 34300 24444 34356
rect 24500 34300 24510 34356
rect 24658 34300 24668 34356
rect 24724 34300 25788 34356
rect 25844 34300 26684 34356
rect 26740 34300 26750 34356
rect 26898 34300 26908 34356
rect 26964 34300 28028 34356
rect 28084 34300 28094 34356
rect 28578 34300 28588 34356
rect 28644 34300 30716 34356
rect 30772 34300 32508 34356
rect 32564 34300 32574 34356
rect 48066 34300 48076 34356
rect 48132 34300 49800 34356
rect 14924 34244 14980 34300
rect 12226 34188 12236 34244
rect 12292 34188 12796 34244
rect 12852 34188 12862 34244
rect 14924 34188 15932 34244
rect 15988 34188 15998 34244
rect 19394 34188 19404 34244
rect 19460 34188 19852 34244
rect 19908 34188 19918 34244
rect 13234 34076 13244 34132
rect 13300 34076 14812 34132
rect 14868 34076 14878 34132
rect 16706 34076 16716 34132
rect 16772 34076 19292 34132
rect 19348 34076 19358 34132
rect 22540 34020 22596 34300
rect 49200 34272 49800 34300
rect 24210 34188 24220 34244
rect 24276 34188 25004 34244
rect 25060 34188 25070 34244
rect 25638 34188 25676 34244
rect 25732 34188 25742 34244
rect 25890 34188 25900 34244
rect 25956 34188 29820 34244
rect 29876 34188 29886 34244
rect 30146 34188 30156 34244
rect 30212 34188 35644 34244
rect 35700 34188 35710 34244
rect 23090 34076 23100 34132
rect 23156 34076 25452 34132
rect 25508 34076 25518 34132
rect 25676 34076 29372 34132
rect 29428 34076 29438 34132
rect 30940 34076 32172 34132
rect 32228 34076 32238 34132
rect 25676 34020 25732 34076
rect 30940 34020 30996 34076
rect 10546 33964 10556 34020
rect 10612 33964 14924 34020
rect 14980 33964 14990 34020
rect 16594 33964 16604 34020
rect 16660 33964 22596 34020
rect 23874 33964 23884 34020
rect 23940 33964 24220 34020
rect 24276 33964 24286 34020
rect 24742 33964 24780 34020
rect 24836 33964 24846 34020
rect 24994 33964 25004 34020
rect 25060 33964 25732 34020
rect 26562 33964 26572 34020
rect 26628 33964 26796 34020
rect 26852 33964 30380 34020
rect 30436 33964 30996 34020
rect 31154 33964 31164 34020
rect 31220 33964 40236 34020
rect 40292 33964 40302 34020
rect 12450 33852 12460 33908
rect 12516 33852 18508 33908
rect 18564 33852 18574 33908
rect 22866 33852 22876 33908
rect 22932 33852 23548 33908
rect 23604 33852 28028 33908
rect 28084 33852 29036 33908
rect 29092 33852 29102 33908
rect 31266 33852 31276 33908
rect 31332 33852 47740 33908
rect 47796 33852 47806 33908
rect 10994 33740 11004 33796
rect 11060 33740 12796 33796
rect 12852 33740 12862 33796
rect 17042 33740 17052 33796
rect 17108 33740 17724 33796
rect 17780 33740 17790 33796
rect 21970 33740 21980 33796
rect 22036 33740 22988 33796
rect 23044 33740 23054 33796
rect 23426 33740 23436 33796
rect 23492 33740 23660 33796
rect 23716 33740 24220 33796
rect 24276 33740 24286 33796
rect 27010 33740 27020 33796
rect 27076 33740 29540 33796
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 29484 33684 29540 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 8306 33628 8316 33684
rect 8372 33628 12572 33684
rect 12628 33628 14700 33684
rect 14756 33628 14766 33684
rect 15092 33628 19404 33684
rect 19460 33628 19470 33684
rect 22204 33628 23548 33684
rect 23604 33628 23614 33684
rect 24770 33628 24780 33684
rect 24836 33628 24892 33684
rect 24948 33628 24958 33684
rect 27122 33628 27132 33684
rect 27188 33628 28924 33684
rect 28980 33628 28990 33684
rect 29474 33628 29484 33684
rect 29540 33628 31164 33684
rect 31220 33628 31230 33684
rect 15092 33572 15148 33628
rect 22204 33572 22260 33628
rect 6626 33516 6636 33572
rect 6692 33516 7980 33572
rect 8036 33516 8046 33572
rect 11106 33516 11116 33572
rect 11172 33516 15148 33572
rect 15810 33516 15820 33572
rect 15876 33516 17276 33572
rect 17332 33516 17342 33572
rect 18358 33516 18396 33572
rect 18452 33516 19852 33572
rect 19908 33516 19918 33572
rect 20850 33516 20860 33572
rect 20916 33516 21308 33572
rect 21364 33516 21374 33572
rect 22194 33516 22204 33572
rect 22260 33516 22270 33572
rect 23762 33516 23772 33572
rect 23828 33516 25004 33572
rect 25060 33516 25070 33572
rect 25666 33516 25676 33572
rect 25732 33516 26908 33572
rect 26964 33516 31276 33572
rect 31332 33516 31342 33572
rect 7980 33348 8036 33516
rect 11330 33404 11340 33460
rect 11396 33404 11676 33460
rect 11732 33404 11742 33460
rect 12114 33404 12124 33460
rect 12180 33404 13580 33460
rect 13636 33404 13646 33460
rect 15474 33404 15484 33460
rect 15540 33404 18732 33460
rect 18788 33404 19740 33460
rect 19796 33404 19806 33460
rect 20066 33404 20076 33460
rect 20132 33404 22316 33460
rect 22372 33404 22382 33460
rect 23202 33404 23212 33460
rect 23268 33404 23660 33460
rect 23716 33404 23726 33460
rect 23958 33404 23996 33460
rect 24052 33404 24062 33460
rect 24882 33404 24892 33460
rect 24948 33404 27468 33460
rect 27524 33404 27534 33460
rect 28130 33404 28140 33460
rect 28196 33404 28812 33460
rect 28868 33404 28878 33460
rect 29698 33404 29708 33460
rect 29764 33404 31948 33460
rect 32004 33404 32732 33460
rect 32788 33404 32798 33460
rect 7980 33292 12348 33348
rect 12404 33292 12414 33348
rect 13010 33292 13020 33348
rect 13076 33292 13086 33348
rect 13346 33292 13356 33348
rect 13412 33292 15036 33348
rect 15092 33292 15102 33348
rect 17042 33292 17052 33348
rect 17108 33292 23884 33348
rect 23940 33292 23950 33348
rect 24518 33292 24556 33348
rect 24612 33292 24622 33348
rect 24882 33292 24892 33348
rect 24948 33292 26908 33348
rect 28690 33292 28700 33348
rect 28756 33292 33852 33348
rect 33908 33292 33918 33348
rect 12534 33180 12572 33236
rect 12628 33180 12638 33236
rect 13020 33124 13076 33292
rect 26852 33236 26908 33292
rect 14578 33180 14588 33236
rect 14644 33180 18788 33236
rect 20178 33180 20188 33236
rect 20244 33180 20636 33236
rect 20692 33180 21868 33236
rect 21924 33180 21934 33236
rect 23650 33180 23660 33236
rect 23716 33180 24780 33236
rect 24836 33180 24846 33236
rect 25414 33180 25452 33236
rect 25508 33180 25518 33236
rect 26852 33180 28700 33236
rect 28756 33180 28766 33236
rect 18732 33124 18788 33180
rect 24780 33124 24836 33180
rect 13020 33068 15820 33124
rect 15876 33068 15886 33124
rect 16258 33068 16268 33124
rect 16324 33068 17612 33124
rect 17668 33068 17678 33124
rect 18722 33068 18732 33124
rect 18788 33068 20860 33124
rect 20916 33068 20926 33124
rect 21522 33068 21532 33124
rect 21588 33068 23324 33124
rect 23380 33068 23548 33124
rect 23604 33068 23614 33124
rect 23762 33068 23772 33124
rect 23828 33068 24108 33124
rect 24164 33068 24174 33124
rect 24780 33068 26012 33124
rect 26068 33068 26078 33124
rect 26450 33068 26460 33124
rect 26516 33068 28252 33124
rect 28308 33068 28318 33124
rect 28466 33068 28476 33124
rect 28532 33068 36988 33124
rect 37044 33068 37054 33124
rect 200 33012 800 33040
rect 200 32956 1820 33012
rect 1876 32956 1886 33012
rect 13010 32956 13020 33012
rect 13076 32956 13468 33012
rect 13524 32956 13534 33012
rect 16118 32956 16156 33012
rect 16212 32956 16222 33012
rect 16370 32956 16380 33012
rect 16436 32956 16474 33012
rect 16594 32956 16604 33012
rect 16660 32956 16716 33012
rect 16772 32956 16782 33012
rect 23426 32956 23436 33012
rect 23492 32956 25564 33012
rect 25620 32956 25630 33012
rect 27458 32956 27468 33012
rect 27524 32956 29260 33012
rect 29316 32956 34412 33012
rect 34468 32956 34478 33012
rect 200 32928 800 32956
rect 16604 32900 16660 32956
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 13570 32844 13580 32900
rect 13636 32844 16660 32900
rect 20188 32844 24556 32900
rect 24612 32844 25228 32900
rect 25284 32844 25294 32900
rect 28354 32844 28364 32900
rect 28420 32844 28476 32900
rect 28532 32844 28542 32900
rect 20188 32788 20244 32844
rect 11890 32732 11900 32788
rect 11956 32732 14924 32788
rect 14980 32732 16828 32788
rect 16884 32732 16894 32788
rect 17378 32732 17388 32788
rect 17444 32732 20244 32788
rect 21298 32732 21308 32788
rect 21364 32732 23548 32788
rect 23604 32732 23614 32788
rect 23846 32732 23884 32788
rect 23940 32732 23950 32788
rect 24882 32732 24892 32788
rect 24948 32732 25676 32788
rect 25732 32732 31052 32788
rect 31108 32732 31118 32788
rect 12226 32620 12236 32676
rect 12292 32620 15596 32676
rect 15652 32620 16716 32676
rect 16772 32620 16782 32676
rect 17266 32620 17276 32676
rect 17332 32620 22036 32676
rect 22502 32620 22540 32676
rect 22596 32620 22606 32676
rect 22866 32620 22876 32676
rect 22932 32620 23436 32676
rect 23492 32620 23502 32676
rect 23958 32620 23996 32676
rect 24052 32620 24668 32676
rect 24724 32620 24734 32676
rect 26002 32620 26012 32676
rect 26068 32620 28700 32676
rect 28756 32620 28766 32676
rect 21980 32564 22036 32620
rect 15362 32508 15372 32564
rect 15428 32508 17388 32564
rect 17444 32508 17454 32564
rect 21970 32508 21980 32564
rect 22036 32508 23772 32564
rect 23828 32508 23838 32564
rect 24994 32508 25004 32564
rect 25060 32508 27244 32564
rect 27300 32508 27310 32564
rect 36082 32508 36092 32564
rect 36148 32508 37996 32564
rect 38052 32508 38062 32564
rect 12002 32396 12012 32452
rect 12068 32396 12236 32452
rect 12292 32396 12302 32452
rect 14018 32396 14028 32452
rect 14084 32396 16380 32452
rect 16436 32396 16446 32452
rect 17714 32396 17724 32452
rect 17780 32396 21308 32452
rect 21364 32396 21374 32452
rect 23762 32396 23772 32452
rect 23828 32396 24332 32452
rect 24388 32396 24398 32452
rect 26534 32396 26572 32452
rect 26628 32396 26638 32452
rect 30146 32396 30156 32452
rect 30212 32396 38668 32452
rect 14466 32284 14476 32340
rect 14532 32284 16828 32340
rect 16884 32284 16894 32340
rect 17042 32284 17052 32340
rect 17108 32284 17164 32340
rect 17220 32284 18508 32340
rect 18564 32284 18574 32340
rect 18732 32284 21532 32340
rect 21588 32284 21598 32340
rect 24210 32284 24220 32340
rect 24276 32284 28476 32340
rect 28532 32284 28542 32340
rect 38612 32284 38668 32396
rect 49200 32340 49800 32368
rect 38724 32284 38734 32340
rect 48066 32284 48076 32340
rect 48132 32284 49800 32340
rect 18732 32228 18788 32284
rect 49200 32256 49800 32284
rect 16146 32172 16156 32228
rect 16212 32172 18788 32228
rect 18844 32172 20748 32228
rect 20804 32172 20814 32228
rect 20962 32172 20972 32228
rect 21028 32172 29708 32228
rect 29764 32172 29774 32228
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 18844 32116 18900 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 15698 32060 15708 32116
rect 15764 32060 16492 32116
rect 16548 32060 18900 32116
rect 19506 32060 19516 32116
rect 19572 32060 19628 32116
rect 19684 32060 19694 32116
rect 20402 32060 20412 32116
rect 20468 32060 21084 32116
rect 21140 32060 21150 32116
rect 21308 32060 26908 32116
rect 21308 32004 21364 32060
rect 12562 31948 12572 32004
rect 12628 31948 16268 32004
rect 16324 31948 16334 32004
rect 16492 31948 17724 32004
rect 17780 31948 17790 32004
rect 18172 31948 18284 32004
rect 18340 31948 18350 32004
rect 19058 31948 19068 32004
rect 19124 31948 19964 32004
rect 20020 31948 20030 32004
rect 20178 31948 20188 32004
rect 20244 31948 20254 32004
rect 20738 31948 20748 32004
rect 20804 31948 21364 32004
rect 22204 31948 22652 32004
rect 22708 31948 22718 32004
rect 16492 31892 16548 31948
rect 18172 31892 18228 31948
rect 20188 31892 20244 31948
rect 22204 31892 22260 31948
rect 10994 31836 11004 31892
rect 11060 31836 16548 31892
rect 16706 31836 16716 31892
rect 16772 31836 17836 31892
rect 17892 31836 17902 31892
rect 18050 31836 18060 31892
rect 18116 31836 18228 31892
rect 18386 31836 18396 31892
rect 18452 31836 18620 31892
rect 18676 31836 19180 31892
rect 19236 31836 19246 31892
rect 19404 31836 21252 31892
rect 21634 31836 21644 31892
rect 21700 31836 22260 31892
rect 22418 31836 22428 31892
rect 22484 31836 22988 31892
rect 23044 31836 23054 31892
rect 25666 31836 25676 31892
rect 25732 31836 25788 31892
rect 25844 31836 25854 31892
rect 19404 31780 19460 31836
rect 10882 31724 10892 31780
rect 10948 31724 16100 31780
rect 16370 31724 16380 31780
rect 16436 31724 18508 31780
rect 18564 31724 18574 31780
rect 18722 31724 18732 31780
rect 18788 31724 19460 31780
rect 200 31584 800 31696
rect 16044 31668 16100 31724
rect 11330 31612 11340 31668
rect 11396 31612 15876 31668
rect 16034 31612 16044 31668
rect 16100 31612 18732 31668
rect 18788 31612 18798 31668
rect 19058 31612 19068 31668
rect 19124 31612 19740 31668
rect 19796 31612 19806 31668
rect 15820 31556 15876 31612
rect 14662 31500 14700 31556
rect 14756 31500 14766 31556
rect 15820 31500 17500 31556
rect 17556 31500 17566 31556
rect 18498 31500 18508 31556
rect 18564 31500 18844 31556
rect 18900 31500 19404 31556
rect 19460 31500 19470 31556
rect 19628 31500 20972 31556
rect 21028 31500 21038 31556
rect 19628 31444 19684 31500
rect 13794 31388 13804 31444
rect 13860 31388 16660 31444
rect 16930 31388 16940 31444
rect 16996 31388 19684 31444
rect 21196 31444 21252 31836
rect 26852 31780 26908 32060
rect 30930 31836 30940 31892
rect 30996 31836 37660 31892
rect 37716 31836 37726 31892
rect 22642 31724 22652 31780
rect 22708 31724 25340 31780
rect 25396 31724 25406 31780
rect 25890 31724 25900 31780
rect 25956 31724 26572 31780
rect 26628 31724 26638 31780
rect 26852 31724 32844 31780
rect 32900 31724 32910 31780
rect 33058 31724 33068 31780
rect 33124 31724 39004 31780
rect 39060 31724 39070 31780
rect 22418 31612 22428 31668
rect 22484 31612 23044 31668
rect 23202 31612 23212 31668
rect 23268 31612 23548 31668
rect 23604 31612 29540 31668
rect 30258 31612 30268 31668
rect 30324 31612 33852 31668
rect 33908 31612 33918 31668
rect 22988 31556 23044 31612
rect 22194 31500 22204 31556
rect 22260 31500 22652 31556
rect 22708 31500 22718 31556
rect 22988 31500 26124 31556
rect 26180 31500 26190 31556
rect 26338 31500 26348 31556
rect 26404 31500 26796 31556
rect 26852 31500 26862 31556
rect 26348 31444 26404 31500
rect 21196 31388 21532 31444
rect 21588 31388 23212 31444
rect 23268 31388 23278 31444
rect 23436 31388 26404 31444
rect 26562 31388 26572 31444
rect 26628 31388 29260 31444
rect 29316 31388 29326 31444
rect 16604 31332 16660 31388
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 9090 31276 9100 31332
rect 9156 31276 16380 31332
rect 16436 31276 16446 31332
rect 16604 31276 17332 31332
rect 17826 31276 17836 31332
rect 17892 31276 19068 31332
rect 19124 31276 19134 31332
rect 21970 31276 21980 31332
rect 22036 31276 23100 31332
rect 23156 31276 23166 31332
rect 17276 31220 17332 31276
rect 23436 31220 23492 31388
rect 29484 31332 29540 31612
rect 24434 31276 24444 31332
rect 24500 31276 26628 31332
rect 29484 31276 32508 31332
rect 32564 31276 32574 31332
rect 14130 31164 14140 31220
rect 14196 31164 14812 31220
rect 14868 31164 14878 31220
rect 15026 31164 15036 31220
rect 15092 31164 16940 31220
rect 16996 31164 17006 31220
rect 17266 31164 17276 31220
rect 17332 31164 18732 31220
rect 18788 31164 18798 31220
rect 19730 31164 19740 31220
rect 19796 31164 23492 31220
rect 19740 31108 19796 31164
rect 26572 31108 26628 31276
rect 26786 31164 26796 31220
rect 26852 31164 34748 31220
rect 34804 31164 34814 31220
rect 19058 31052 19068 31108
rect 19124 31052 19796 31108
rect 21186 31052 21196 31108
rect 21252 31052 23996 31108
rect 24052 31052 24062 31108
rect 26114 31052 26124 31108
rect 26180 31052 26190 31108
rect 26572 31052 37436 31108
rect 37492 31052 37502 31108
rect 26124 30996 26180 31052
rect 49200 30996 49800 31024
rect 9426 30940 9436 30996
rect 9492 30940 15596 30996
rect 15652 30940 17164 30996
rect 17220 30940 17230 30996
rect 17938 30940 17948 30996
rect 18004 30940 18172 30996
rect 18228 30940 20524 30996
rect 20580 30940 20590 30996
rect 21186 30940 21196 30996
rect 21252 30940 26068 30996
rect 26124 30940 28924 30996
rect 28980 30940 28990 30996
rect 29250 30940 29260 30996
rect 29316 30940 36652 30996
rect 36708 30940 36718 30996
rect 48066 30940 48076 30996
rect 48132 30940 49800 30996
rect 26012 30884 26068 30940
rect 49200 30912 49800 30940
rect 12114 30828 12124 30884
rect 12180 30828 17724 30884
rect 17780 30828 19068 30884
rect 19124 30828 19134 30884
rect 22418 30828 22428 30884
rect 22484 30828 24444 30884
rect 24500 30828 24510 30884
rect 26012 30828 26124 30884
rect 26180 30828 36764 30884
rect 36820 30828 36830 30884
rect 14802 30716 14812 30772
rect 14868 30716 19068 30772
rect 19124 30716 19134 30772
rect 19730 30716 19740 30772
rect 19796 30716 20524 30772
rect 20580 30716 20860 30772
rect 20916 30716 20926 30772
rect 21634 30716 21644 30772
rect 21700 30716 22988 30772
rect 23044 30716 23054 30772
rect 10658 30604 10668 30660
rect 10724 30604 15820 30660
rect 15876 30604 16604 30660
rect 16660 30604 16670 30660
rect 16818 30604 16828 30660
rect 16884 30604 20188 30660
rect 20244 30604 20254 30660
rect 20402 30604 20412 30660
rect 20468 30604 23884 30660
rect 23940 30604 23950 30660
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 7522 30492 7532 30548
rect 7588 30492 18060 30548
rect 18116 30492 19068 30548
rect 19124 30492 19628 30548
rect 19684 30492 19694 30548
rect 20188 30492 20748 30548
rect 20804 30492 26236 30548
rect 26292 30492 26302 30548
rect 20188 30436 20244 30492
rect 17154 30380 17164 30436
rect 17220 30380 20244 30436
rect 20402 30380 20412 30436
rect 20468 30380 20860 30436
rect 20916 30380 21644 30436
rect 21700 30380 21710 30436
rect 24434 30380 24444 30436
rect 24500 30380 28252 30436
rect 28308 30380 28318 30436
rect 17266 30268 17276 30324
rect 17332 30268 17836 30324
rect 17892 30268 18396 30324
rect 18452 30268 18462 30324
rect 19404 30212 19460 30380
rect 19618 30268 19628 30324
rect 19684 30268 20748 30324
rect 20804 30268 20814 30324
rect 23986 30268 23996 30324
rect 24052 30268 25116 30324
rect 25172 30268 25182 30324
rect 9986 30156 9996 30212
rect 10052 30156 16044 30212
rect 16100 30156 16110 30212
rect 19170 30156 19180 30212
rect 19236 30156 19460 30212
rect 19516 30156 20860 30212
rect 20916 30156 20926 30212
rect 22642 30156 22652 30212
rect 22708 30156 23436 30212
rect 23492 30156 23884 30212
rect 23940 30156 23950 30212
rect 26002 30156 26012 30212
rect 26068 30156 26796 30212
rect 26852 30156 30828 30212
rect 30884 30156 30894 30212
rect 19516 30100 19572 30156
rect 8866 30044 8876 30100
rect 8932 30044 15260 30100
rect 15316 30044 15326 30100
rect 15484 30044 19572 30100
rect 19842 30044 19852 30100
rect 19908 30044 21140 30100
rect 21298 30044 21308 30100
rect 21364 30044 28588 30100
rect 28644 30044 28654 30100
rect 29362 30044 29372 30100
rect 29428 30044 29932 30100
rect 29988 30044 29998 30100
rect 15484 29988 15540 30044
rect 21084 29988 21140 30044
rect 15138 29932 15148 29988
rect 15204 29932 15540 29988
rect 18732 29932 20300 29988
rect 20356 29932 20366 29988
rect 21084 29932 24780 29988
rect 24836 29932 34972 29988
rect 35028 29932 35038 29988
rect 18732 29876 18788 29932
rect 13906 29820 13916 29876
rect 13972 29820 18732 29876
rect 18788 29820 18798 29876
rect 20514 29820 20524 29876
rect 20580 29820 20590 29876
rect 20850 29820 20860 29876
rect 20916 29820 21196 29876
rect 21252 29820 27804 29876
rect 27860 29820 27870 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 9202 29708 9212 29764
rect 9268 29708 19180 29764
rect 19236 29708 19404 29764
rect 19460 29708 19470 29764
rect 200 29652 800 29680
rect 20524 29652 20580 29820
rect 20962 29708 20972 29764
rect 21028 29708 34524 29764
rect 34580 29708 34590 29764
rect 200 29596 1820 29652
rect 1876 29596 1886 29652
rect 18610 29596 18620 29652
rect 18676 29596 19404 29652
rect 19460 29596 19740 29652
rect 19796 29596 19806 29652
rect 20524 29596 20860 29652
rect 20916 29596 21364 29652
rect 23090 29596 23100 29652
rect 23156 29596 36540 29652
rect 36596 29596 36606 29652
rect 200 29568 800 29596
rect 21308 29540 21364 29596
rect 5506 29484 5516 29540
rect 5572 29484 21084 29540
rect 21140 29484 21150 29540
rect 21308 29484 30604 29540
rect 30660 29484 30670 29540
rect 15922 29372 15932 29428
rect 15988 29372 21196 29428
rect 21252 29372 21262 29428
rect 16594 29260 16604 29316
rect 16660 29260 20860 29316
rect 20916 29260 20926 29316
rect 21568 29260 21644 29316
rect 21700 29260 35084 29316
rect 35140 29260 35150 29316
rect 19394 29148 19404 29204
rect 19460 29148 22876 29204
rect 22932 29148 22942 29204
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 49200 28980 49800 29008
rect 48066 28924 48076 28980
rect 48132 28924 49800 28980
rect 49200 28896 49800 28924
rect 21904 28700 21980 28756
rect 22036 28700 22540 28756
rect 22596 28700 22606 28756
rect 22978 28700 22988 28756
rect 23044 28700 23212 28756
rect 23268 28700 32620 28756
rect 32676 28700 32686 28756
rect 8978 28476 8988 28532
rect 9044 28476 18620 28532
rect 18676 28476 19628 28532
rect 19684 28476 19694 28532
rect 24770 28476 24780 28532
rect 24836 28476 30604 28532
rect 30660 28476 30670 28532
rect 200 28308 800 28336
rect 200 28252 1820 28308
rect 1876 28252 1886 28308
rect 26852 28252 36876 28308
rect 36932 28252 36942 28308
rect 200 28224 800 28252
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 26852 28196 26908 28252
rect 26226 28140 26236 28196
rect 26292 28140 26908 28196
rect 28578 28140 28588 28196
rect 28644 28140 31948 28196
rect 32004 28140 32014 28196
rect 19058 28028 19068 28084
rect 19124 28028 32956 28084
rect 33012 28028 33022 28084
rect 6738 27916 6748 27972
rect 6804 27916 26460 27972
rect 26516 27916 26526 27972
rect 6290 27804 6300 27860
rect 6356 27804 21532 27860
rect 21588 27804 21598 27860
rect 20514 27580 20524 27636
rect 20580 27580 35980 27636
rect 36036 27580 36046 27636
rect 15474 27468 15484 27524
rect 15540 27468 30044 27524
rect 30100 27468 30110 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 10882 27356 10892 27412
rect 10948 27356 20412 27412
rect 20468 27356 20478 27412
rect 19618 27244 19628 27300
rect 19684 27244 36988 27300
rect 37044 27244 37054 27300
rect 18050 27132 18060 27188
rect 18116 27132 30268 27188
rect 30324 27132 30334 27188
rect 49200 26964 49800 26992
rect 48076 26908 49800 26964
rect 48076 26852 48132 26908
rect 49200 26880 49800 26908
rect 8306 26796 8316 26852
rect 8372 26796 22540 26852
rect 22596 26796 22606 26852
rect 33842 26796 33852 26852
rect 33908 26796 37212 26852
rect 37268 26796 37278 26852
rect 48066 26796 48076 26852
rect 48132 26796 48142 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 16370 26460 16380 26516
rect 16436 26460 30940 26516
rect 30996 26460 31006 26516
rect 16706 26348 16716 26404
rect 16772 26348 28588 26404
rect 28644 26348 28654 26404
rect 200 26292 800 26320
rect 200 26236 1820 26292
rect 1876 26236 1886 26292
rect 12338 26236 12348 26292
rect 12404 26236 29932 26292
rect 29988 26236 29998 26292
rect 200 26208 800 26236
rect 6514 26124 6524 26180
rect 6580 26124 22764 26180
rect 22820 26124 22830 26180
rect 16594 25900 16604 25956
rect 16660 25900 31276 25956
rect 31332 25900 31342 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 14690 25788 14700 25844
rect 14756 25788 31164 25844
rect 31220 25788 31230 25844
rect 49200 25536 49800 25648
rect 26898 25116 26908 25172
rect 26964 25116 28476 25172
rect 28532 25116 36540 25172
rect 36596 25116 36606 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 13122 24892 13132 24948
rect 13188 24892 32844 24948
rect 32900 24892 32910 24948
rect 8530 24780 8540 24836
rect 8596 24780 26124 24836
rect 26180 24780 26190 24836
rect 18386 24668 18396 24724
rect 18452 24668 30268 24724
rect 30324 24668 30334 24724
rect 20132 24556 21756 24612
rect 21812 24556 21822 24612
rect 22418 24556 22428 24612
rect 22484 24556 35756 24612
rect 35812 24556 35822 24612
rect 20132 24500 20188 24556
rect 4162 24444 4172 24500
rect 4228 24444 19628 24500
rect 19684 24444 20188 24500
rect 200 24276 800 24304
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 200 24220 1820 24276
rect 1876 24220 1886 24276
rect 12338 24220 12348 24276
rect 12404 24220 33180 24276
rect 33236 24220 33246 24276
rect 200 24192 800 24220
rect 7746 24108 7756 24164
rect 7812 24108 26908 24164
rect 26964 24108 26974 24164
rect 19058 23996 19068 24052
rect 19124 23996 32060 24052
rect 32116 23996 32126 24052
rect 12898 23660 12908 23716
rect 12964 23660 22988 23716
rect 23044 23660 23054 23716
rect 49200 23604 49800 23632
rect 48066 23548 48076 23604
rect 48132 23548 49800 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 49200 23520 49800 23548
rect 1922 23324 1932 23380
rect 1988 23324 17836 23380
rect 17892 23324 17902 23380
rect 7298 23212 7308 23268
rect 7364 23212 28140 23268
rect 28196 23212 40460 23268
rect 40516 23212 40526 23268
rect 200 22932 800 22960
rect 200 22876 2044 22932
rect 2100 22876 2110 22932
rect 200 22848 800 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 11666 21756 11676 21812
rect 11732 21756 40348 21812
rect 40404 21756 40414 21812
rect 12786 21644 12796 21700
rect 12852 21644 36428 21700
rect 36484 21644 36494 21700
rect 49200 21588 49800 21616
rect 13570 21532 13580 21588
rect 13636 21532 36316 21588
rect 36372 21532 36382 21588
rect 48066 21532 48076 21588
rect 48132 21532 49800 21588
rect 49200 21504 49800 21532
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 200 20916 800 20944
rect 200 20860 1820 20916
rect 1876 20860 1886 20916
rect 200 20832 800 20860
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 49200 20160 49800 20272
rect 2930 20076 2940 20132
rect 2996 20076 33292 20132
rect 33348 20076 33358 20132
rect 11554 19964 11564 20020
rect 11620 19964 33628 20020
rect 33684 19964 33694 20020
rect 22754 19852 22764 19908
rect 22820 19852 40012 19908
rect 40068 19852 40078 19908
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 200 18900 800 18928
rect 200 18844 1820 18900
rect 1876 18844 1886 18900
rect 200 18816 800 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 48066 18508 48076 18564
rect 48132 18508 48142 18564
rect 6962 18396 6972 18452
rect 7028 18396 42028 18452
rect 42084 18396 42094 18452
rect 3938 18284 3948 18340
rect 4004 18284 31948 18340
rect 32004 18284 32014 18340
rect 48076 18228 48132 18508
rect 49200 18228 49800 18256
rect 3490 18172 3500 18228
rect 3556 18172 22652 18228
rect 22708 18172 22718 18228
rect 48076 18172 49800 18228
rect 49200 18144 49800 18172
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 200 17556 800 17584
rect 200 17500 1820 17556
rect 1876 17500 1886 17556
rect 200 17472 800 17500
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 49200 16884 49800 16912
rect 48066 16828 48076 16884
rect 48132 16828 49800 16884
rect 49200 16800 49800 16828
rect 16146 16716 16156 16772
rect 16212 16716 36092 16772
rect 36148 16716 36158 16772
rect 20962 16604 20972 16660
rect 21028 16604 38780 16660
rect 38836 16604 38846 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 15026 16380 15036 16436
rect 15092 16380 24108 16436
rect 24164 16380 24174 16436
rect 22978 16268 22988 16324
rect 23044 16268 39452 16324
rect 39508 16268 39518 16324
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 200 15540 800 15568
rect 200 15484 1820 15540
rect 1876 15484 1886 15540
rect 200 15456 800 15484
rect 6626 15036 6636 15092
rect 6692 15036 35644 15092
rect 35700 15036 35710 15092
rect 4834 14924 4844 14980
rect 4900 14924 26012 14980
rect 26068 14924 26078 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 10546 14812 10556 14868
rect 10612 14812 21980 14868
rect 22036 14812 23436 14868
rect 23492 14812 23502 14868
rect 49200 14784 49800 14896
rect 200 14196 800 14224
rect 200 14140 1820 14196
rect 1876 14140 1886 14196
rect 200 14112 800 14140
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 22642 13244 22652 13300
rect 22708 13244 34188 13300
rect 34244 13244 34254 13300
rect 23426 13132 23436 13188
rect 23492 13132 40348 13188
rect 40404 13132 40414 13188
rect 49200 12852 49800 12880
rect 48066 12796 48076 12852
rect 48132 12796 49800 12852
rect 49200 12768 49800 12796
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 200 12096 800 12208
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 6626 11676 6636 11732
rect 6692 11676 23772 11732
rect 23828 11676 23838 11732
rect 10658 11564 10668 11620
rect 10724 11564 26572 11620
rect 26628 11564 26638 11620
rect 49200 11508 49800 11536
rect 19394 11452 19404 11508
rect 19460 11452 29372 11508
rect 29428 11452 29438 11508
rect 48066 11452 48076 11508
rect 48132 11452 49800 11508
rect 49200 11424 49800 11452
rect 19618 11340 19628 11396
rect 19684 11340 38668 11396
rect 38724 11340 38734 11396
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 200 10164 800 10192
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 200 10108 1820 10164
rect 1876 10108 1886 10164
rect 200 10080 800 10108
rect 7410 9772 7420 9828
rect 7476 9772 9100 9828
rect 9156 9772 9166 9828
rect 9090 9548 9100 9604
rect 9156 9548 9548 9604
rect 9604 9548 12684 9604
rect 12740 9548 12750 9604
rect 49200 9492 49800 9520
rect 48066 9436 48076 9492
rect 48132 9436 49800 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 49200 9408 49800 9436
rect 200 8820 800 8848
rect 200 8764 1820 8820
rect 1876 8764 1886 8820
rect 200 8736 800 8764
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 49200 7476 49800 7504
rect 48066 7420 48076 7476
rect 48132 7420 49800 7476
rect 49200 7392 49800 7420
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 200 6804 800 6832
rect 200 6748 1820 6804
rect 1876 6748 1886 6804
rect 200 6720 800 6748
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 49200 6132 49800 6160
rect 48066 6076 48076 6132
rect 48132 6076 49800 6132
rect 49200 6048 49800 6076
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 200 4704 800 4816
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 49200 4032 49800 4144
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 3042 3612 3052 3668
rect 3108 3612 4284 3668
rect 4340 3612 8764 3668
rect 8820 3612 8830 3668
rect 1362 3500 1372 3556
rect 1428 3500 2156 3556
rect 2212 3500 2222 3556
rect 200 3444 800 3472
rect 200 3388 1820 3444
rect 1876 3388 1886 3444
rect 36418 3388 36428 3444
rect 36484 3388 36988 3444
rect 37044 3388 37548 3444
rect 37604 3388 37614 3444
rect 47506 3388 47516 3444
rect 47572 3388 48076 3444
rect 48132 3388 49084 3444
rect 49140 3388 49150 3444
rect 200 3360 800 3388
rect 4722 3276 4732 3332
rect 4788 3276 5740 3332
rect 5796 3276 5806 3332
rect 28242 3276 28252 3332
rect 28308 3276 29260 3332
rect 29316 3276 29326 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 18 2268 28 2324
rect 84 2268 2492 2324
rect 2548 2268 2558 2324
rect 49200 2100 49800 2128
rect 48178 2044 48188 2100
rect 48244 2044 49800 2100
rect 49200 2016 49800 2044
rect 200 1344 800 1456
rect 49200 756 49800 784
rect 47170 700 47180 756
rect 47236 700 49800 756
rect 49200 672 49800 700
<< via3 >>
rect 34748 49868 34804 49924
rect 11676 49756 11732 49812
rect 25788 49644 25844 49700
rect 18956 49532 19012 49588
rect 9548 49420 9604 49476
rect 26012 49420 26068 49476
rect 30492 49420 30548 49476
rect 26348 49308 26404 49364
rect 26012 49196 26068 49252
rect 26796 49196 26852 49252
rect 11564 49084 11620 49140
rect 27804 48860 27860 48916
rect 25788 48636 25844 48692
rect 16604 48524 16660 48580
rect 16940 48524 16996 48580
rect 29036 48524 29092 48580
rect 26796 48412 26852 48468
rect 27356 48412 27412 48468
rect 36316 48300 36372 48356
rect 7980 48188 8036 48244
rect 30380 48188 30436 48244
rect 8372 47964 8428 48020
rect 11340 47964 11396 48020
rect 14028 47964 14084 48020
rect 34300 47964 34356 48020
rect 7868 47852 7924 47908
rect 15596 47852 15652 47908
rect 29596 47852 29652 47908
rect 8316 47628 8372 47684
rect 14924 47628 14980 47684
rect 16716 47516 16772 47572
rect 25452 47516 25508 47572
rect 36316 47404 36372 47460
rect 27356 47292 27412 47348
rect 27580 47292 27636 47348
rect 29148 47180 29204 47236
rect 33292 47180 33348 47236
rect 8540 47068 8596 47124
rect 10332 47068 10388 47124
rect 27468 47068 27524 47124
rect 8316 46956 8372 47012
rect 24556 46956 24612 47012
rect 17948 46620 18004 46676
rect 29932 46620 29988 46676
rect 29260 46508 29316 46564
rect 10780 46396 10836 46452
rect 27692 46396 27748 46452
rect 31052 46284 31108 46340
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 33628 46172 33684 46228
rect 11788 46060 11844 46116
rect 13244 46060 13300 46116
rect 17724 45948 17780 46004
rect 27692 45948 27748 46004
rect 24556 45836 24612 45892
rect 35868 45836 35924 45892
rect 13468 45612 13524 45668
rect 28364 45612 28420 45668
rect 31500 45612 31556 45668
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 29484 45500 29540 45556
rect 29820 45500 29876 45556
rect 30156 45500 30212 45556
rect 11452 45388 11508 45444
rect 30268 45388 30324 45444
rect 7868 45164 7924 45220
rect 10108 45164 10164 45220
rect 7980 45052 8036 45108
rect 11340 45052 11396 45108
rect 11788 45052 11844 45108
rect 19628 45052 19684 45108
rect 28140 45052 28196 45108
rect 29708 45052 29764 45108
rect 33404 45052 33460 45108
rect 36876 44940 36932 44996
rect 10556 44828 10612 44884
rect 12348 44828 12404 44884
rect 29484 44716 29540 44772
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 30268 44604 30324 44660
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 31388 44492 31444 44548
rect 31612 44492 31668 44548
rect 4172 44380 4228 44436
rect 14812 44380 14868 44436
rect 40460 44380 40516 44436
rect 11564 44268 11620 44324
rect 14700 44268 14756 44324
rect 10332 44156 10388 44212
rect 25116 44156 25172 44212
rect 8988 44044 9044 44100
rect 10780 44044 10836 44100
rect 27692 44044 27748 44100
rect 29708 44044 29764 44100
rect 34412 43932 34468 43988
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 29372 43820 29428 43876
rect 10668 43708 10724 43764
rect 11900 43708 11956 43764
rect 12460 43708 12516 43764
rect 25900 43708 25956 43764
rect 33516 43708 33572 43764
rect 10780 43596 10836 43652
rect 11788 43596 11844 43652
rect 14812 43596 14868 43652
rect 30268 43596 30324 43652
rect 30604 43596 30660 43652
rect 36764 43596 36820 43652
rect 11228 43484 11284 43540
rect 12460 43484 12516 43540
rect 24108 43484 24164 43540
rect 31276 43484 31332 43540
rect 35756 43484 35812 43540
rect 18060 43372 18116 43428
rect 21532 43372 21588 43428
rect 29036 43372 29092 43428
rect 30380 43372 30436 43428
rect 29708 43260 29764 43316
rect 29932 43260 29988 43316
rect 34188 43260 34244 43316
rect 37436 43260 37492 43316
rect 40348 43260 40404 43316
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 31836 43148 31892 43204
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 26908 43036 26964 43092
rect 36204 43036 36260 43092
rect 18060 42924 18116 42980
rect 20972 42812 21028 42868
rect 28588 42812 28644 42868
rect 31164 42700 31220 42756
rect 8204 42588 8260 42644
rect 9100 42588 9156 42644
rect 23772 42588 23828 42644
rect 30604 42588 30660 42644
rect 30940 42588 30996 42644
rect 31612 42588 31668 42644
rect 37436 42588 37492 42644
rect 9324 42476 9380 42532
rect 32956 42476 33012 42532
rect 34860 42476 34916 42532
rect 39452 42476 39508 42532
rect 14700 42364 14756 42420
rect 18508 42364 18564 42420
rect 20860 42364 20916 42420
rect 29036 42364 29092 42420
rect 30716 42364 30772 42420
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 33404 42364 33460 42420
rect 35756 42364 35812 42420
rect 9772 42252 9828 42308
rect 36204 42252 36260 42308
rect 6972 42028 7028 42084
rect 8540 42028 8596 42084
rect 10892 42028 10948 42084
rect 18172 42140 18228 42196
rect 26908 42140 26964 42196
rect 28700 42140 28756 42196
rect 31164 42140 31220 42196
rect 29036 42028 29092 42084
rect 29484 42028 29540 42084
rect 31276 42028 31332 42084
rect 33068 42140 33124 42196
rect 31948 42028 32004 42084
rect 34748 42028 34804 42084
rect 39004 42028 39060 42084
rect 6412 41916 6468 41972
rect 29820 41916 29876 41972
rect 30044 41916 30100 41972
rect 35644 41916 35700 41972
rect 35980 41916 36036 41972
rect 36988 41916 37044 41972
rect 3500 41804 3556 41860
rect 4956 41804 5012 41860
rect 8316 41804 8372 41860
rect 23548 41804 23604 41860
rect 32172 41804 32228 41860
rect 6636 41692 6692 41748
rect 7308 41692 7364 41748
rect 19516 41692 19572 41748
rect 30380 41692 30436 41748
rect 33516 41692 33572 41748
rect 34972 41692 35028 41748
rect 4844 41580 4900 41636
rect 10780 41580 10836 41636
rect 34076 41580 34132 41636
rect 35644 41580 35700 41636
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 6636 41468 6692 41524
rect 30156 41468 30212 41524
rect 35868 41468 35924 41524
rect 7980 41356 8036 41412
rect 8652 41356 8708 41412
rect 8876 41356 8932 41412
rect 25004 41356 25060 41412
rect 9548 41244 9604 41300
rect 29260 41244 29316 41300
rect 29596 41244 29652 41300
rect 31500 41244 31556 41300
rect 31836 41244 31892 41300
rect 35644 41244 35700 41300
rect 8316 41132 8372 41188
rect 23548 41132 23604 41188
rect 32620 41132 32676 41188
rect 33404 41132 33460 41188
rect 3500 41020 3556 41076
rect 4844 41020 4900 41076
rect 7308 41020 7364 41076
rect 20188 41020 20244 41076
rect 23660 41020 23716 41076
rect 28476 41020 28532 41076
rect 29708 41020 29764 41076
rect 28812 40908 28868 40964
rect 32396 40908 32452 40964
rect 32732 40908 32788 40964
rect 33180 40908 33236 40964
rect 36428 40908 36484 40964
rect 37436 40908 37492 40964
rect 39004 40908 39060 40964
rect 8876 40796 8932 40852
rect 10444 40796 10500 40852
rect 37100 40796 37156 40852
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 7980 40684 8036 40740
rect 16716 40684 16772 40740
rect 30380 40684 30436 40740
rect 33740 40684 33796 40740
rect 29596 40572 29652 40628
rect 31612 40572 31668 40628
rect 13356 40460 13412 40516
rect 15932 40460 15988 40516
rect 20188 40460 20244 40516
rect 29484 40460 29540 40516
rect 31836 40460 31892 40516
rect 32508 40460 32564 40516
rect 9660 40348 9716 40404
rect 12012 40348 12068 40404
rect 15708 40348 15764 40404
rect 18284 40348 18340 40404
rect 24444 40348 24500 40404
rect 30940 40348 30996 40404
rect 33068 40348 33124 40404
rect 33964 40348 34020 40404
rect 36204 40348 36260 40404
rect 38780 40348 38836 40404
rect 11004 40236 11060 40292
rect 13580 40236 13636 40292
rect 29372 40236 29428 40292
rect 29596 40236 29652 40292
rect 30268 40236 30324 40292
rect 33740 40236 33796 40292
rect 34412 40236 34468 40292
rect 8652 40124 8708 40180
rect 29260 40124 29316 40180
rect 32284 40124 32340 40180
rect 32732 40124 32788 40180
rect 7868 40012 7924 40068
rect 26796 40012 26852 40068
rect 31500 40012 31556 40068
rect 34412 40012 34468 40068
rect 34860 40012 34916 40068
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 15036 39900 15092 39956
rect 21756 39900 21812 39956
rect 29932 39900 29988 39956
rect 33292 39900 33348 39956
rect 33740 39900 33796 39956
rect 30044 39788 30100 39844
rect 30604 39788 30660 39844
rect 30828 39788 30884 39844
rect 7420 39676 7476 39732
rect 21644 39676 21700 39732
rect 30268 39676 30324 39732
rect 31164 39676 31220 39732
rect 9772 39564 9828 39620
rect 15036 39564 15092 39620
rect 24780 39564 24836 39620
rect 30716 39564 30772 39620
rect 33292 39564 33348 39620
rect 33628 39564 33684 39620
rect 13580 39452 13636 39508
rect 18732 39452 18788 39508
rect 9436 39340 9492 39396
rect 29260 39340 29316 39396
rect 30268 39340 30324 39396
rect 7868 39228 7924 39284
rect 15372 39228 15428 39284
rect 27916 39228 27972 39284
rect 33516 39228 33572 39284
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 9772 39116 9828 39172
rect 31836 39116 31892 39172
rect 33292 39116 33348 39172
rect 10556 39004 10612 39060
rect 10108 38892 10164 38948
rect 17164 38892 17220 38948
rect 27804 38892 27860 38948
rect 28812 38892 28868 38948
rect 30156 38892 30212 38948
rect 30380 38892 30436 38948
rect 31052 38892 31108 38948
rect 32956 38892 33012 38948
rect 8428 38780 8484 38836
rect 18844 38780 18900 38836
rect 19628 38780 19684 38836
rect 30044 38780 30100 38836
rect 33852 38780 33908 38836
rect 38668 38780 38724 38836
rect 7420 38668 7476 38724
rect 10556 38668 10612 38724
rect 13244 38668 13300 38724
rect 21868 38668 21924 38724
rect 24556 38668 24612 38724
rect 28028 38668 28084 38724
rect 15372 38556 15428 38612
rect 16156 38556 16212 38612
rect 19516 38556 19572 38612
rect 32508 38668 32564 38724
rect 28700 38556 28756 38612
rect 30268 38556 30324 38612
rect 34300 38556 34356 38612
rect 36540 38556 36596 38612
rect 30380 38444 30436 38500
rect 35868 38444 35924 38500
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 12012 38332 12068 38388
rect 27580 38332 27636 38388
rect 31612 38332 31668 38388
rect 30828 38220 30884 38276
rect 31500 38220 31556 38276
rect 10780 38108 10836 38164
rect 13468 38108 13524 38164
rect 31724 38108 31780 38164
rect 34300 38108 34356 38164
rect 36540 38108 36596 38164
rect 19068 37996 19124 38052
rect 28700 37996 28756 38052
rect 29036 37996 29092 38052
rect 35868 37996 35924 38052
rect 36764 37996 36820 38052
rect 10332 37884 10388 37940
rect 10556 37884 10612 37940
rect 34860 37884 34916 37940
rect 11900 37772 11956 37828
rect 13244 37772 13300 37828
rect 13468 37772 13524 37828
rect 15036 37772 15092 37828
rect 28700 37772 28756 37828
rect 30268 37772 30324 37828
rect 33180 37772 33236 37828
rect 37100 37772 37156 37828
rect 18956 37660 19012 37716
rect 33964 37660 34020 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 12012 37548 12068 37604
rect 29484 37548 29540 37604
rect 29932 37548 29988 37604
rect 11564 37436 11620 37492
rect 34076 37436 34132 37492
rect 34636 37436 34692 37492
rect 8764 37324 8820 37380
rect 8988 37324 9044 37380
rect 9996 37324 10052 37380
rect 10556 37324 10612 37380
rect 13244 37324 13300 37380
rect 28588 37324 28644 37380
rect 28812 37324 28868 37380
rect 30492 37324 30548 37380
rect 34748 37324 34804 37380
rect 16380 37212 16436 37268
rect 20188 37212 20244 37268
rect 21868 37212 21924 37268
rect 28028 37212 28084 37268
rect 28364 37212 28420 37268
rect 21756 37100 21812 37156
rect 26236 37100 26292 37156
rect 31612 37100 31668 37156
rect 36540 37100 36596 37156
rect 9324 36988 9380 37044
rect 10556 36988 10612 37044
rect 16380 36988 16436 37044
rect 23100 36988 23156 37044
rect 30380 36988 30436 37044
rect 30604 36988 30660 37044
rect 33404 36988 33460 37044
rect 36204 36988 36260 37044
rect 4844 36876 4900 36932
rect 9660 36876 9716 36932
rect 21868 36876 21924 36932
rect 27356 36876 27412 36932
rect 32620 36876 32676 36932
rect 33852 36876 33908 36932
rect 34300 36876 34356 36932
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 28476 36764 28532 36820
rect 12572 36652 12628 36708
rect 32284 36652 32340 36708
rect 38780 36652 38836 36708
rect 6412 36540 6468 36596
rect 8428 36540 8484 36596
rect 17836 36540 17892 36596
rect 21756 36540 21812 36596
rect 23772 36540 23828 36596
rect 14028 36428 14084 36484
rect 35868 36428 35924 36484
rect 17724 36316 17780 36372
rect 22988 36316 23044 36372
rect 26796 36316 26852 36372
rect 6748 36204 6804 36260
rect 8204 36204 8260 36260
rect 12124 36204 12180 36260
rect 28812 36204 28868 36260
rect 30044 36204 30100 36260
rect 30716 36204 30772 36260
rect 31836 36204 31892 36260
rect 8652 36092 8708 36148
rect 13692 36092 13748 36148
rect 25900 36092 25956 36148
rect 32956 36092 33012 36148
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 9996 35980 10052 36036
rect 10444 35980 10500 36036
rect 12124 35980 12180 36036
rect 31388 35980 31444 36036
rect 11788 35868 11844 35924
rect 27692 35868 27748 35924
rect 28476 35868 28532 35924
rect 29148 35868 29204 35924
rect 15036 35756 15092 35812
rect 23100 35756 23156 35812
rect 24780 35756 24836 35812
rect 28588 35756 28644 35812
rect 31724 35644 31780 35700
rect 7308 35532 7364 35588
rect 9100 35532 9156 35588
rect 18508 35532 18564 35588
rect 25676 35532 25732 35588
rect 27356 35532 27412 35588
rect 27580 35532 27636 35588
rect 20188 35420 20244 35476
rect 26124 35420 26180 35476
rect 32732 35420 32788 35476
rect 6524 35308 6580 35364
rect 25116 35308 25172 35364
rect 29596 35308 29652 35364
rect 30828 35308 30884 35364
rect 32172 35308 32228 35364
rect 33068 35308 33124 35364
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 13692 35196 13748 35252
rect 14924 35196 14980 35252
rect 27916 35196 27972 35252
rect 28252 35196 28308 35252
rect 33964 35196 34020 35252
rect 27020 35084 27076 35140
rect 31276 35084 31332 35140
rect 21644 34860 21700 34916
rect 14700 34748 14756 34804
rect 16380 34748 16436 34804
rect 32396 34748 32452 34804
rect 11228 34636 11284 34692
rect 25004 34636 25060 34692
rect 16492 34524 16548 34580
rect 25900 34524 25956 34580
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 15092 34300 15148 34356
rect 20860 34300 20916 34356
rect 24444 34300 24500 34356
rect 25788 34300 25844 34356
rect 26684 34300 26740 34356
rect 28588 34300 28644 34356
rect 32508 34300 32564 34356
rect 12236 34188 12292 34244
rect 12796 34188 12852 34244
rect 14812 34076 14868 34132
rect 25676 34188 25732 34244
rect 25900 34188 25956 34244
rect 35644 34188 35700 34244
rect 23884 33964 23940 34020
rect 24780 33964 24836 34020
rect 26572 33964 26628 34020
rect 30380 33964 30436 34020
rect 31164 33964 31220 34020
rect 27020 33740 27076 33796
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 23548 33628 23604 33684
rect 24892 33628 24948 33684
rect 18396 33516 18452 33572
rect 25676 33516 25732 33572
rect 11340 33404 11396 33460
rect 23996 33404 24052 33460
rect 29708 33404 29764 33460
rect 24556 33292 24612 33348
rect 24892 33292 24948 33348
rect 28700 33292 28756 33348
rect 12572 33180 12628 33236
rect 23660 33180 23716 33236
rect 25452 33180 25508 33236
rect 21532 33068 21588 33124
rect 28252 33068 28308 33124
rect 13468 32956 13524 33012
rect 16156 32956 16212 33012
rect 16380 32956 16436 33012
rect 16604 32956 16660 33012
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 24556 32844 24612 32900
rect 28476 32844 28532 32900
rect 23884 32732 23940 32788
rect 22540 32620 22596 32676
rect 23996 32620 24052 32676
rect 28700 32620 28756 32676
rect 23772 32508 23828 32564
rect 12012 32396 12068 32452
rect 16380 32396 16436 32452
rect 26572 32396 26628 32452
rect 30156 32396 30212 32452
rect 17164 32284 17220 32340
rect 38668 32284 38724 32340
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 16492 32060 16548 32116
rect 19628 32060 19684 32116
rect 19068 31948 19124 32004
rect 11004 31836 11060 31892
rect 22428 31836 22484 31892
rect 25788 31836 25844 31892
rect 18732 31724 18788 31780
rect 14700 31500 14756 31556
rect 18844 31500 18900 31556
rect 30940 31836 30996 31892
rect 33068 31724 33124 31780
rect 39004 31724 39060 31780
rect 33852 31612 33908 31668
rect 22652 31500 22708 31556
rect 29260 31388 29316 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 24444 31276 24500 31332
rect 18732 31164 18788 31220
rect 21196 31052 21252 31108
rect 37436 31052 37492 31108
rect 9436 30940 9492 30996
rect 28924 30940 28980 30996
rect 29260 30940 29316 30996
rect 12124 30828 12180 30884
rect 19068 30828 19124 30884
rect 22428 30828 22484 30884
rect 20524 30716 20580 30772
rect 20860 30716 20916 30772
rect 20188 30604 20244 30660
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 26236 30492 26292 30548
rect 20412 30380 20468 30436
rect 21644 30380 21700 30436
rect 18396 30268 18452 30324
rect 19628 30268 19684 30324
rect 9996 30156 10052 30212
rect 23436 30156 23492 30212
rect 26012 30156 26068 30212
rect 26796 30156 26852 30212
rect 30828 30156 30884 30212
rect 8876 30044 8932 30100
rect 28588 30044 28644 30100
rect 29372 30044 29428 30100
rect 29932 30044 29988 30100
rect 34972 29932 35028 29988
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 19180 29708 19236 29764
rect 19404 29708 19460 29764
rect 15932 29372 15988 29428
rect 21196 29372 21252 29428
rect 21644 29260 21700 29316
rect 19404 29148 19460 29204
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 21980 28700 22036 28756
rect 22540 28700 22596 28756
rect 8988 28476 9044 28532
rect 18620 28476 18676 28532
rect 19628 28476 19684 28532
rect 24780 28476 24836 28532
rect 30604 28476 30660 28532
rect 36876 28252 36932 28308
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 26236 28140 26292 28196
rect 31948 28140 32004 28196
rect 19068 28028 19124 28084
rect 6748 27916 6804 27972
rect 20524 27580 20580 27636
rect 35980 27580 36036 27636
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 10892 27356 10948 27412
rect 19628 27244 19684 27300
rect 36988 27244 37044 27300
rect 18060 27132 18116 27188
rect 30268 27132 30324 27188
rect 8316 26796 8372 26852
rect 22540 26796 22596 26852
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 16380 26460 16436 26516
rect 30940 26460 30996 26516
rect 6524 26124 6580 26180
rect 16604 25900 16660 25956
rect 31276 25900 31332 25956
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 14700 25788 14756 25844
rect 31164 25788 31220 25844
rect 26908 25116 26964 25172
rect 28476 25116 28532 25172
rect 36540 25116 36596 25172
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 32844 24892 32900 24948
rect 8540 24780 8596 24836
rect 26124 24780 26180 24836
rect 35756 24556 35812 24612
rect 4172 24444 4228 24500
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 12348 24220 12404 24276
rect 33180 24220 33236 24276
rect 26908 24108 26964 24164
rect 22988 23660 23044 23716
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 17836 23324 17892 23380
rect 28140 23212 28196 23268
rect 40460 23212 40516 23268
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 12796 21644 12852 21700
rect 36428 21644 36484 21700
rect 13580 21532 13636 21588
rect 36316 21532 36372 21588
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 33292 20076 33348 20132
rect 11564 19964 11620 20020
rect 33628 19964 33684 20020
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 6972 18396 7028 18452
rect 3500 18172 3556 18228
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 20972 16604 21028 16660
rect 38780 16604 38836 16660
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 24108 16380 24164 16436
rect 22988 16268 23044 16324
rect 39452 16268 39508 16324
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4844 14924 4900 14980
rect 26012 14924 26068 14980
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 10556 14812 10612 14868
rect 21980 14812 22036 14868
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 22652 13244 22708 13300
rect 34188 13244 34244 13300
rect 40348 13132 40404 13188
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 6636 11676 6692 11732
rect 10668 11564 10724 11620
rect 26572 11564 26628 11620
rect 29372 11452 29428 11508
rect 38668 11340 38724 11396
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 7420 9772 7476 9828
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 34748 49924 34804 49934
rect 11676 49812 11732 49822
rect 9548 49476 9604 49486
rect 7980 48244 8036 48254
rect 7868 47908 7924 47918
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 7868 45220 7924 47852
rect 7868 45154 7924 45164
rect 7980 45108 8036 48188
rect 8372 48020 8428 48030
rect 8428 47964 8596 48020
rect 8372 47954 8428 47964
rect 8316 47684 8372 47694
rect 8316 47012 8372 47628
rect 8540 47124 8596 47964
rect 8540 47058 8596 47068
rect 8316 46946 8372 46956
rect 7980 45042 8036 45052
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4172 44436 4228 44446
rect 3500 41860 3556 41870
rect 3500 41076 3556 41804
rect 3500 18228 3556 41020
rect 4172 24500 4228 44380
rect 4172 24434 4228 24444
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 8988 44100 9044 44110
rect 8204 42644 8260 42654
rect 6972 42084 7028 42094
rect 6412 41972 6468 41982
rect 4956 41860 5012 41870
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4844 41636 4900 41646
rect 4844 41076 4900 41580
rect 4844 41010 4900 41020
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4956 38668 5012 41804
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 3500 18162 3556 18172
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4844 38612 5012 38668
rect 4844 36932 4900 38612
rect 4844 14980 4900 36876
rect 6412 36596 6468 41916
rect 6412 36530 6468 36540
rect 6636 41748 6692 41758
rect 6636 41524 6692 41692
rect 6524 35364 6580 35374
rect 6524 26180 6580 35308
rect 6524 26114 6580 26124
rect 4844 14914 4900 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 6636 11732 6692 41468
rect 6748 36260 6804 36270
rect 6748 27972 6804 36204
rect 6748 27906 6804 27916
rect 6972 18452 7028 42028
rect 7308 41748 7364 41758
rect 7308 41076 7364 41692
rect 7308 35588 7364 41020
rect 7980 41412 8036 41422
rect 7980 40740 8036 41356
rect 7980 40674 8036 40684
rect 7868 40068 7924 40078
rect 7308 35522 7364 35532
rect 7420 39732 7476 39742
rect 7420 38724 7476 39676
rect 7868 39284 7924 40012
rect 7868 39218 7924 39228
rect 6972 18386 7028 18396
rect 6636 11666 6692 11676
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 7420 9828 7476 38668
rect 8204 36260 8260 42588
rect 8540 42084 8596 42094
rect 8204 36194 8260 36204
rect 8316 41860 8372 41870
rect 8316 41188 8372 41804
rect 8316 26852 8372 41132
rect 8428 38836 8484 38846
rect 8428 36596 8484 38780
rect 8428 36530 8484 36540
rect 8316 26786 8372 26796
rect 8540 24836 8596 42028
rect 8652 41412 8708 41422
rect 8876 41412 8932 41422
rect 8708 41356 8820 41412
rect 8652 41346 8708 41356
rect 8652 40180 8708 40190
rect 8652 36148 8708 40124
rect 8764 37380 8820 41356
rect 8876 40852 8932 41356
rect 8876 40786 8932 40796
rect 8988 38668 9044 44044
rect 8764 37314 8820 37324
rect 8876 38612 9044 38668
rect 9100 42644 9156 42654
rect 8652 36082 8708 36092
rect 8876 30100 8932 38612
rect 8876 30034 8932 30044
rect 8988 37380 9044 37390
rect 8988 28532 9044 37324
rect 9100 35588 9156 42588
rect 9324 42532 9380 42542
rect 9324 37044 9380 42476
rect 9548 41300 9604 49420
rect 11564 49140 11620 49150
rect 11340 49084 11564 49140
rect 11340 48020 11396 49084
rect 11564 49074 11620 49084
rect 11340 47954 11396 47964
rect 10332 47124 10388 47134
rect 10108 45220 10164 45230
rect 9548 41234 9604 41244
rect 9772 42308 9828 42318
rect 9660 40404 9716 40414
rect 9324 36978 9380 36988
rect 9436 39396 9492 39406
rect 9100 35522 9156 35532
rect 9436 30996 9492 39340
rect 9660 36932 9716 40348
rect 9772 39620 9828 42252
rect 9772 39172 9828 39564
rect 9772 39106 9828 39116
rect 10108 38948 10164 45164
rect 10108 38882 10164 38892
rect 10332 44212 10388 47068
rect 10780 46452 10836 46462
rect 10332 37940 10388 44156
rect 10556 44884 10612 44894
rect 10332 37874 10388 37884
rect 10444 40852 10500 40862
rect 9660 36866 9716 36876
rect 9996 37380 10052 37390
rect 9436 30930 9492 30940
rect 9996 36036 10052 37324
rect 9996 30212 10052 35980
rect 10444 36036 10500 40796
rect 10556 39060 10612 44828
rect 10780 44100 10836 46396
rect 11452 45444 11508 45454
rect 10556 38724 10612 39004
rect 10556 38658 10612 38668
rect 10668 43764 10724 43774
rect 10556 37940 10612 37950
rect 10556 37380 10612 37884
rect 10556 37314 10612 37324
rect 10444 35970 10500 35980
rect 10556 37044 10612 37054
rect 9996 30146 10052 30156
rect 8988 28466 9044 28476
rect 8540 24770 8596 24780
rect 10556 14868 10612 36988
rect 10556 14802 10612 14812
rect 10668 11620 10724 43708
rect 10780 43652 10836 44044
rect 10780 43586 10836 43596
rect 11340 45108 11396 45118
rect 11228 43540 11284 43550
rect 10892 42084 10948 42094
rect 10780 41636 10836 41646
rect 10780 38164 10836 41580
rect 10780 38098 10836 38108
rect 10892 27412 10948 42028
rect 11004 40292 11060 40302
rect 11004 31892 11060 40236
rect 11228 34692 11284 43484
rect 11228 34626 11284 34636
rect 11340 33460 11396 45052
rect 11340 33394 11396 33404
rect 11004 31826 11060 31836
rect 10892 27346 10948 27356
rect 11452 26908 11508 45388
rect 11564 44324 11620 44334
rect 11564 37492 11620 44268
rect 11676 43876 11732 49756
rect 25788 49700 25844 49710
rect 18956 49588 19012 49598
rect 16604 48580 16660 48590
rect 16940 48580 16996 48590
rect 16660 48524 16940 48580
rect 16604 48514 16660 48524
rect 16940 48514 16996 48524
rect 14028 48020 14084 48030
rect 11788 46116 11844 46126
rect 11788 45108 11844 46060
rect 11788 45042 11844 45052
rect 13244 46116 13300 46126
rect 12348 44884 12404 44894
rect 11676 43820 11956 43876
rect 11900 43764 11956 43820
rect 11900 43698 11956 43708
rect 11564 37426 11620 37436
rect 11788 43652 11844 43662
rect 11788 35924 11844 43596
rect 12012 40404 12068 40414
rect 12012 38668 12068 40348
rect 11900 38612 12292 38668
rect 11900 37828 11956 38612
rect 11900 37762 11956 37772
rect 12012 38388 12068 38398
rect 11788 35858 11844 35868
rect 12012 37604 12068 38332
rect 12012 32452 12068 37548
rect 12012 32386 12068 32396
rect 12124 36260 12180 36270
rect 12124 36036 12180 36204
rect 12124 30884 12180 35980
rect 12236 34244 12292 38612
rect 12236 34178 12292 34188
rect 12124 30818 12180 30828
rect 11452 26852 11620 26908
rect 11564 20020 11620 26852
rect 12348 24276 12404 44828
rect 12460 43764 12516 43774
rect 12460 43540 12516 43708
rect 12460 43474 12516 43484
rect 13244 38724 13300 46060
rect 13468 45668 13524 45678
rect 13468 43708 13524 45612
rect 13356 43652 13524 43708
rect 13356 40516 13412 43652
rect 13356 40450 13412 40460
rect 13244 38658 13300 38668
rect 13580 40292 13636 40302
rect 13580 39508 13636 40236
rect 13468 38164 13524 38174
rect 13244 37828 13300 37838
rect 13244 37380 13300 37772
rect 13244 37314 13300 37324
rect 13468 37828 13524 38108
rect 12572 36708 12628 36718
rect 12572 33236 12628 36652
rect 12572 33170 12628 33180
rect 12796 34244 12852 34254
rect 12348 24210 12404 24220
rect 12796 21700 12852 34188
rect 13468 33012 13524 37772
rect 13468 32946 13524 32956
rect 12796 21634 12852 21644
rect 13580 21588 13636 39452
rect 14028 36484 14084 47964
rect 15596 47908 15652 47918
rect 15652 47852 15764 47908
rect 15596 47842 15652 47852
rect 14924 47684 14980 47694
rect 14812 44436 14868 44446
rect 14700 44324 14756 44334
rect 14700 42420 14756 44268
rect 14700 42354 14756 42364
rect 14812 43652 14868 44380
rect 14028 36418 14084 36428
rect 13692 36148 13748 36158
rect 13692 35252 13748 36092
rect 13692 35186 13748 35196
rect 14700 34804 14756 34814
rect 14700 31556 14756 34748
rect 14812 34468 14868 43596
rect 14924 35252 14980 47628
rect 15708 40404 15764 47852
rect 16716 47572 16772 47582
rect 16716 40740 16772 47516
rect 17948 46676 18004 46686
rect 15708 40338 15764 40348
rect 15932 40516 15988 40526
rect 15036 39956 15092 39966
rect 15036 39620 15092 39900
rect 15036 37828 15092 39564
rect 15372 39284 15428 39294
rect 15372 38612 15428 39228
rect 15372 38546 15428 38556
rect 15036 35812 15092 37772
rect 15036 35746 15092 35756
rect 14924 35186 14980 35196
rect 14812 34412 15092 34468
rect 14812 34132 14868 34412
rect 15036 34366 15092 34412
rect 15036 34356 15148 34366
rect 15036 34300 15092 34356
rect 15092 34290 15148 34300
rect 14812 34066 14868 34076
rect 14700 25844 14756 31500
rect 15932 29428 15988 40460
rect 16716 38668 16772 40684
rect 17724 46004 17780 46014
rect 16156 38612 16212 38622
rect 16156 33012 16212 38556
rect 16604 38612 16772 38668
rect 17164 38948 17220 38958
rect 16380 37268 16436 37278
rect 16380 37044 16436 37212
rect 16380 36978 16436 36988
rect 16156 32946 16212 32956
rect 16380 34804 16436 34814
rect 16380 33012 16436 34748
rect 15932 29362 15988 29372
rect 16380 32452 16436 32956
rect 16380 26516 16436 32396
rect 16492 34580 16548 34590
rect 16492 32116 16548 34524
rect 16492 32050 16548 32060
rect 16604 33012 16660 38612
rect 16380 26450 16436 26460
rect 16604 25956 16660 32956
rect 17164 32340 17220 38892
rect 17724 36372 17780 45948
rect 17948 38668 18004 46620
rect 17724 36306 17780 36316
rect 17836 38612 18004 38668
rect 18060 43428 18116 43438
rect 18060 42980 18116 43372
rect 17836 36596 17892 38612
rect 17164 32274 17220 32284
rect 16604 25890 16660 25900
rect 14700 25778 14756 25788
rect 17836 23380 17892 36540
rect 18060 27188 18116 42924
rect 18508 42420 18564 42430
rect 18172 42196 18228 42206
rect 18228 42140 18340 42196
rect 18172 42130 18228 42140
rect 18284 40404 18340 42140
rect 18284 40338 18340 40348
rect 18508 35588 18564 42364
rect 18732 39508 18788 39518
rect 18732 38668 18788 39452
rect 18508 35522 18564 35532
rect 18620 38612 18788 38668
rect 18844 38836 18900 38846
rect 18396 33572 18452 33582
rect 18396 30324 18452 33516
rect 18396 30258 18452 30268
rect 18620 28532 18676 38612
rect 18732 31780 18788 31790
rect 18732 31220 18788 31724
rect 18844 31556 18900 38780
rect 18956 37716 19012 49532
rect 25788 48692 25844 49644
rect 26012 49476 26068 49486
rect 26012 49252 26068 49420
rect 30492 49476 30548 49486
rect 26348 49364 26404 49374
rect 26404 49308 26852 49364
rect 26348 49298 26404 49308
rect 26012 49186 26068 49196
rect 26796 49252 26852 49308
rect 26796 49186 26852 49196
rect 25788 48626 25844 48636
rect 27804 48916 27860 48926
rect 26796 48468 26852 48478
rect 25452 47572 25508 47582
rect 24556 47012 24612 47022
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19628 45108 19684 45118
rect 19516 41748 19572 41758
rect 19516 38612 19572 41692
rect 19516 38546 19572 38556
rect 19628 38836 19684 45052
rect 18956 37650 19012 37660
rect 19068 38052 19124 38062
rect 19068 35308 19124 37996
rect 19068 35252 19236 35308
rect 18844 31490 18900 31500
rect 19068 32004 19124 32014
rect 18732 31154 18788 31164
rect 18620 28466 18676 28476
rect 19068 30884 19124 31948
rect 19068 28084 19124 30828
rect 19180 29764 19236 35252
rect 19628 32116 19684 38780
rect 19628 30324 19684 32060
rect 19628 30258 19684 30268
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 24556 45892 24612 46956
rect 24108 43540 24164 43550
rect 21532 43428 21588 43438
rect 20972 42868 21028 42878
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 20860 42420 20916 42430
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 20188 41076 20244 41086
rect 20188 40516 20244 41020
rect 20188 40450 20244 40460
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 20188 37268 20244 37278
rect 20188 35476 20244 37212
rect 20188 35410 20244 35420
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 20860 34356 20916 42364
rect 20524 30772 20580 30782
rect 20188 30660 20244 30670
rect 20188 30436 20244 30604
rect 20412 30436 20468 30446
rect 20188 30380 20412 30436
rect 20412 30370 20468 30380
rect 19180 29698 19236 29708
rect 19404 29764 19460 29774
rect 19404 29204 19460 29708
rect 19404 29138 19460 29148
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19068 28018 19124 28028
rect 19628 28532 19684 28542
rect 19628 27300 19684 28476
rect 19628 27234 19684 27244
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 18060 27122 18116 27132
rect 17836 23314 17892 23324
rect 19808 26684 20128 28196
rect 20524 27636 20580 30716
rect 20860 30772 20916 34300
rect 20860 30706 20916 30716
rect 20524 27570 20580 27580
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 13580 21522 13636 21532
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 11564 19954 11620 19964
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 10668 11554 10724 11564
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 20972 16660 21028 42812
rect 21532 33124 21588 43372
rect 23772 42644 23828 42654
rect 23548 41860 23604 41870
rect 23548 41188 23604 41804
rect 21756 39956 21812 39966
rect 21644 39732 21700 39742
rect 21644 34916 21700 39676
rect 21756 37156 21812 39900
rect 21868 38724 21924 38734
rect 21868 38612 23044 38668
rect 21756 36596 21812 37100
rect 21868 37268 21924 37278
rect 21868 36932 21924 37212
rect 21868 36866 21924 36876
rect 21756 36530 21812 36540
rect 21644 34850 21700 34860
rect 22988 36372 23044 38612
rect 21532 33058 21588 33068
rect 22540 32676 22596 32686
rect 22428 31892 22484 31902
rect 21196 31108 21252 31118
rect 21196 29428 21252 31052
rect 22428 30884 22484 31836
rect 21196 29362 21252 29372
rect 21644 30436 21700 30446
rect 21644 29316 21700 30380
rect 21644 29250 21700 29260
rect 20972 16594 21028 16604
rect 21980 28756 22036 28766
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 21980 14868 22036 28700
rect 22428 26908 22484 30828
rect 22540 28756 22596 32620
rect 22540 28690 22596 28700
rect 22652 31556 22708 31566
rect 22428 26852 22596 26908
rect 22540 26786 22596 26796
rect 21980 14802 22036 14812
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 22652 13300 22708 31500
rect 22988 23716 23044 36316
rect 23100 37044 23156 37054
rect 23100 35812 23156 36988
rect 23100 35746 23156 35756
rect 23548 33684 23604 41132
rect 23436 33628 23548 33684
rect 23436 30212 23492 33628
rect 23548 33618 23604 33628
rect 23660 41076 23716 41086
rect 23660 33236 23716 41020
rect 23660 33170 23716 33180
rect 23772 36596 23828 42588
rect 23772 32564 23828 36540
rect 23884 34020 23940 34030
rect 23884 32788 23940 33964
rect 23884 32722 23940 32732
rect 23996 33460 24052 33470
rect 23996 32676 24052 33404
rect 23996 32610 24052 32620
rect 23772 32498 23828 32508
rect 23436 30146 23492 30156
rect 22988 16324 23044 23660
rect 24108 16436 24164 43484
rect 24444 40404 24500 40414
rect 24444 34356 24500 40348
rect 24556 38724 24612 45836
rect 25116 44212 25172 44222
rect 25004 41412 25060 41422
rect 24556 38658 24612 38668
rect 24780 39620 24836 39630
rect 24780 35812 24836 39564
rect 24780 35746 24836 35756
rect 25004 34692 25060 41356
rect 25116 35364 25172 44156
rect 25116 35298 25172 35308
rect 25004 34626 25060 34636
rect 24444 31332 24500 34300
rect 24780 34020 24836 34030
rect 24556 33348 24612 33358
rect 24556 32900 24612 33292
rect 24556 32834 24612 32844
rect 24444 31266 24500 31276
rect 24780 28532 24836 33964
rect 24892 33684 24948 33694
rect 24892 33348 24948 33628
rect 24892 33282 24948 33292
rect 25452 33236 25508 47516
rect 25900 43764 25956 43774
rect 25900 36148 25956 43708
rect 26796 40068 26852 48412
rect 27356 48468 27412 48478
rect 27356 47348 27412 48412
rect 27580 47348 27636 47358
rect 27356 47282 27412 47292
rect 27468 47292 27580 47348
rect 27468 47124 27524 47292
rect 27580 47282 27636 47292
rect 27468 47058 27524 47068
rect 27692 46452 27748 46462
rect 27692 46004 27748 46396
rect 27692 45938 27748 45948
rect 27692 44100 27748 44110
rect 26908 43092 26964 43102
rect 26908 42196 26964 43036
rect 26908 42130 26964 42140
rect 26684 40012 26796 40068
rect 25900 36082 25956 36092
rect 26236 37156 26292 37166
rect 25676 35588 25732 35598
rect 25676 34244 25732 35532
rect 26124 35476 26180 35486
rect 25900 34580 25956 34590
rect 25676 33572 25732 34188
rect 25676 33506 25732 33516
rect 25788 34356 25844 34366
rect 25452 33170 25508 33180
rect 25788 31892 25844 34300
rect 25900 34244 25956 34524
rect 25900 34178 25956 34188
rect 25788 31826 25844 31836
rect 24780 28466 24836 28476
rect 26012 30212 26068 30222
rect 24108 16370 24164 16380
rect 22988 16258 23044 16268
rect 26012 14980 26068 30156
rect 26124 24836 26180 35420
rect 26236 30548 26292 37100
rect 26684 34356 26740 40012
rect 26796 40002 26852 40012
rect 27580 38388 27636 38398
rect 27356 36932 27412 36942
rect 26684 34290 26740 34300
rect 26796 36372 26852 36382
rect 26236 28196 26292 30492
rect 26236 28130 26292 28140
rect 26572 34020 26628 34030
rect 26572 32452 26628 33964
rect 26124 24770 26180 24780
rect 26012 14914 26068 14924
rect 22652 13234 22708 13244
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 7420 9762 7476 9772
rect 19808 11004 20128 12516
rect 26572 11620 26628 32396
rect 26796 30212 26852 36316
rect 27356 35588 27412 36876
rect 27356 35522 27412 35532
rect 27580 35588 27636 38332
rect 27692 35924 27748 44044
rect 27804 38948 27860 48860
rect 29036 48580 29092 48590
rect 28364 45668 28420 45678
rect 28140 45108 28196 45118
rect 27804 38882 27860 38892
rect 27916 39284 27972 39294
rect 27692 35858 27748 35868
rect 27580 35522 27636 35532
rect 27916 35252 27972 39228
rect 28028 38724 28084 38734
rect 28028 37268 28084 38668
rect 28028 37202 28084 37212
rect 27916 35186 27972 35196
rect 27020 35140 27076 35150
rect 27020 33796 27076 35084
rect 27020 33730 27076 33740
rect 26796 30146 26852 30156
rect 26908 25172 26964 25182
rect 26908 24164 26964 25116
rect 26908 24098 26964 24108
rect 28140 23268 28196 45052
rect 28364 37268 28420 45612
rect 29036 43428 29092 48524
rect 30380 48244 30436 48254
rect 29596 47908 29652 47918
rect 28588 42868 28644 42878
rect 28252 35252 28308 35262
rect 28252 33124 28308 35196
rect 28252 33058 28308 33068
rect 28364 26908 28420 37212
rect 28476 41076 28532 41086
rect 28476 36820 28532 41020
rect 28588 37380 28644 42812
rect 29036 42420 29092 43372
rect 28924 42364 29036 42420
rect 28700 42196 28756 42206
rect 28700 38612 28756 42140
rect 28812 40964 28868 40974
rect 28812 38948 28868 40908
rect 28812 38882 28868 38892
rect 28700 38546 28756 38556
rect 28700 38052 28756 38062
rect 28756 37996 28868 38052
rect 28700 37986 28756 37996
rect 28588 37314 28644 37324
rect 28700 37828 28756 37838
rect 28476 36754 28532 36764
rect 28476 35924 28532 35934
rect 28476 32900 28532 35868
rect 28476 32834 28532 32844
rect 28588 35812 28644 35822
rect 28588 34356 28644 35756
rect 28588 30100 28644 34300
rect 28700 33348 28756 37772
rect 28812 37380 28868 37996
rect 28812 36260 28868 37324
rect 28812 36194 28868 36204
rect 28700 32676 28756 33292
rect 28700 32610 28756 32620
rect 28924 30996 28980 42364
rect 29036 42354 29092 42364
rect 29148 47236 29204 47246
rect 29036 42084 29092 42094
rect 29036 38052 29092 42028
rect 29036 37986 29092 37996
rect 29148 35924 29204 47180
rect 29260 46564 29316 46574
rect 29260 41300 29316 46508
rect 29484 45556 29540 45566
rect 29484 44772 29540 45500
rect 29260 41234 29316 41244
rect 29372 43876 29428 43886
rect 29372 40292 29428 43820
rect 29484 42084 29540 44716
rect 29484 42018 29540 42028
rect 29596 41300 29652 47852
rect 29932 46676 29988 46686
rect 29820 45556 29876 45566
rect 29708 45108 29764 45118
rect 29708 44100 29764 45052
rect 29708 44034 29764 44044
rect 29596 41234 29652 41244
rect 29708 43316 29764 43326
rect 29708 41076 29764 43260
rect 29820 41972 29876 45500
rect 29932 45556 29988 46620
rect 30156 45556 30212 45566
rect 29932 45500 30156 45556
rect 29932 43316 29988 45500
rect 30156 45490 30212 45500
rect 30268 45444 30324 45454
rect 30268 44660 30324 45388
rect 30268 43652 30324 44604
rect 30268 43586 30324 43596
rect 29932 43250 29988 43260
rect 30380 43428 30436 48188
rect 29820 41906 29876 41916
rect 30044 41972 30100 41982
rect 29708 41010 29764 41020
rect 29596 40628 29652 40638
rect 29652 40572 29764 40628
rect 29596 40562 29652 40572
rect 29372 40226 29428 40236
rect 29484 40516 29540 40526
rect 29260 40180 29316 40190
rect 29260 39396 29316 40124
rect 29260 39330 29316 39340
rect 29484 37604 29540 40460
rect 29484 37538 29540 37548
rect 29596 40292 29652 40302
rect 29148 35858 29204 35868
rect 29596 35364 29652 40236
rect 29596 35298 29652 35308
rect 29708 33460 29764 40572
rect 29708 33394 29764 33404
rect 29932 39956 29988 39966
rect 29932 37604 29988 39900
rect 30044 39844 30100 41916
rect 30380 41748 30436 43372
rect 30380 41682 30436 41692
rect 30044 39778 30100 39788
rect 30156 41524 30212 41534
rect 30156 38948 30212 41468
rect 30380 40740 30436 40750
rect 30268 40292 30324 40302
rect 30268 39732 30324 40236
rect 30268 39666 30324 39676
rect 28924 30930 28980 30940
rect 29260 31444 29316 31454
rect 29260 30996 29316 31388
rect 29260 30930 29316 30940
rect 28588 30034 28644 30044
rect 29372 30100 29428 30110
rect 28364 26852 28532 26908
rect 28476 25172 28532 26852
rect 28476 25106 28532 25116
rect 28140 23202 28196 23212
rect 26572 11554 26628 11564
rect 29372 11508 29428 30044
rect 29932 30100 29988 37548
rect 30044 38836 30100 38846
rect 30044 36260 30100 38780
rect 30044 36194 30100 36204
rect 30156 32452 30212 38892
rect 30268 39396 30324 39406
rect 30268 38612 30324 39340
rect 30380 38948 30436 40684
rect 30380 38882 30436 38892
rect 30268 38546 30324 38556
rect 30380 38500 30436 38510
rect 30156 32386 30212 32396
rect 30268 37828 30324 37838
rect 29932 30034 29988 30044
rect 30268 27188 30324 37772
rect 30380 37044 30436 38444
rect 30492 37380 30548 49420
rect 34300 48020 34356 48030
rect 33292 47236 33348 47246
rect 31052 46340 31108 46350
rect 30604 43652 30660 43662
rect 30604 42644 30660 43596
rect 30940 42644 30996 42654
rect 30604 42578 30660 42588
rect 30716 42588 30940 42644
rect 30716 42420 30772 42588
rect 30940 42578 30996 42588
rect 30716 42354 30772 42364
rect 30940 40404 30996 40414
rect 30492 37314 30548 37324
rect 30604 39844 30660 39854
rect 30380 34020 30436 36988
rect 30380 33954 30436 33964
rect 30604 37044 30660 39788
rect 30828 39844 30884 39854
rect 30604 28532 30660 36988
rect 30716 39620 30772 39630
rect 30716 36260 30772 39564
rect 30828 38276 30884 39788
rect 30828 38210 30884 38220
rect 30716 36194 30772 36204
rect 30828 35364 30884 35374
rect 30828 30212 30884 35308
rect 30828 30146 30884 30156
rect 30940 31892 30996 40348
rect 31052 38948 31108 46284
rect 31500 45668 31556 45678
rect 31388 44548 31444 44558
rect 31276 43540 31332 43550
rect 31164 42756 31220 42766
rect 31164 42196 31220 42700
rect 31164 42130 31220 42140
rect 31276 42084 31332 43484
rect 31052 38882 31108 38892
rect 31164 39732 31220 39742
rect 30604 28466 30660 28476
rect 30268 27122 30324 27132
rect 30940 26516 30996 31836
rect 30940 26450 30996 26460
rect 31164 34020 31220 39676
rect 31164 25844 31220 33964
rect 31276 35140 31332 42028
rect 31388 36036 31444 44492
rect 31500 44548 31556 45612
rect 31612 44548 31668 44558
rect 31500 44492 31612 44548
rect 31500 41300 31556 44492
rect 31612 44482 31668 44492
rect 31836 43204 31892 43214
rect 31500 41234 31556 41244
rect 31612 42644 31668 42654
rect 31612 40628 31668 42588
rect 31500 40068 31556 40078
rect 31500 38276 31556 40012
rect 31500 38210 31556 38220
rect 31612 38388 31668 40572
rect 31836 41300 31892 43148
rect 32956 42532 33012 42542
rect 31836 40516 31892 41244
rect 31836 40450 31892 40460
rect 31948 42084 32004 42094
rect 31612 37156 31668 38332
rect 31836 39172 31892 39182
rect 31612 37090 31668 37100
rect 31724 38164 31780 38174
rect 31388 35970 31444 35980
rect 31724 35700 31780 38108
rect 31836 36260 31892 39116
rect 31836 36194 31892 36204
rect 31724 35634 31780 35644
rect 31276 25956 31332 35084
rect 31948 28196 32004 42028
rect 32172 41860 32228 41870
rect 32172 41188 32228 41804
rect 32620 41188 32676 41198
rect 32172 41132 32620 41188
rect 32172 35364 32228 41132
rect 32620 41122 32676 41132
rect 32396 40964 32452 40974
rect 32396 40628 32452 40908
rect 32732 40964 32788 40974
rect 32396 40572 32564 40628
rect 32284 40180 32340 40190
rect 32284 36708 32340 40124
rect 32284 36642 32340 36652
rect 32172 35298 32228 35308
rect 32396 34804 32452 40572
rect 32508 40516 32564 40572
rect 32508 40450 32564 40460
rect 32732 40404 32788 40908
rect 32620 40348 32788 40404
rect 32396 34738 32452 34748
rect 32508 38724 32564 38734
rect 32508 34356 32564 38668
rect 32620 36932 32676 40348
rect 32620 36866 32676 36876
rect 32732 40180 32788 40190
rect 32732 35476 32788 40124
rect 32956 39172 33012 42476
rect 33068 42196 33124 42206
rect 33068 40404 33124 42140
rect 33068 40338 33124 40348
rect 33180 40964 33236 40974
rect 32732 35410 32788 35420
rect 32844 39116 33012 39172
rect 32508 34290 32564 34300
rect 31948 28130 32004 28140
rect 31276 25890 31332 25900
rect 31164 25778 31220 25788
rect 32844 24948 32900 39116
rect 32956 38948 33012 38958
rect 32956 36148 33012 38892
rect 33180 38668 33236 40908
rect 33292 39956 33348 47180
rect 33628 46228 33684 46238
rect 33404 45108 33460 45118
rect 33404 42420 33460 45052
rect 33404 42354 33460 42364
rect 33516 43764 33572 43774
rect 33516 41748 33572 43708
rect 33516 41682 33572 41692
rect 33292 39890 33348 39900
rect 33404 41188 33460 41198
rect 33292 39620 33348 39630
rect 33292 39172 33348 39564
rect 33292 39106 33348 39116
rect 33180 38612 33348 38668
rect 32956 36082 33012 36092
rect 33180 37828 33236 37838
rect 33068 35364 33124 35374
rect 33068 31780 33124 35308
rect 33068 31714 33124 31724
rect 32844 24882 32900 24892
rect 33180 24276 33236 37772
rect 33180 24210 33236 24220
rect 33292 20132 33348 38612
rect 33404 37044 33460 41132
rect 33628 39620 33684 46172
rect 34188 43316 34244 43326
rect 34076 41636 34132 41646
rect 33740 40740 33796 40750
rect 33796 40684 33908 40740
rect 33740 40674 33796 40684
rect 33740 40292 33796 40302
rect 33740 39956 33796 40236
rect 33740 39890 33796 39900
rect 33628 39554 33684 39564
rect 33404 36978 33460 36988
rect 33516 39284 33572 39294
rect 33516 35308 33572 39228
rect 33852 38836 33908 40684
rect 33852 38770 33908 38780
rect 33964 40404 34020 40414
rect 33964 37716 34020 40348
rect 33852 36932 33908 36942
rect 33516 35252 33684 35308
rect 33292 20066 33348 20076
rect 33628 20020 33684 35252
rect 33852 31668 33908 36876
rect 33964 35252 34020 37660
rect 34076 37492 34132 41580
rect 34076 37426 34132 37436
rect 33964 35186 34020 35196
rect 33852 31602 33908 31612
rect 33628 19954 33684 19964
rect 34188 13300 34244 43260
rect 34300 38948 34356 47964
rect 34412 43988 34468 43998
rect 34412 40292 34468 43932
rect 34748 42084 34804 49868
rect 36316 48356 36372 48366
rect 36316 47460 36372 48300
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35868 45892 35924 45902
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 34748 42018 34804 42028
rect 34860 42532 34916 42542
rect 34860 41860 34916 42476
rect 34412 40068 34468 40236
rect 34412 40002 34468 40012
rect 34748 41804 34916 41860
rect 34300 38892 34692 38948
rect 34300 38612 34356 38622
rect 34300 38164 34356 38556
rect 34300 36932 34356 38108
rect 34636 37492 34692 38892
rect 34636 37426 34692 37436
rect 34748 37380 34804 41804
rect 34972 41748 35028 41758
rect 34860 40068 34916 40078
rect 34860 37940 34916 40012
rect 34860 37874 34916 37884
rect 34748 37314 34804 37324
rect 34300 36866 34356 36876
rect 34972 29988 35028 41692
rect 34972 29922 35028 29932
rect 35168 41580 35488 43092
rect 35756 43540 35812 43550
rect 35756 42420 35812 43484
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35644 41972 35700 41982
rect 35644 41636 35700 41916
rect 35644 41570 35700 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35644 41300 35700 41310
rect 35644 34244 35700 41244
rect 35644 34178 35700 34188
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 34188 13234 34244 13244
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35756 24612 35812 42364
rect 35868 41524 35924 45836
rect 36204 43092 36260 43102
rect 36204 42308 36260 43036
rect 36204 42242 36260 42252
rect 35868 38500 35924 41468
rect 35868 38434 35924 38444
rect 35980 41972 36036 41982
rect 35868 38052 35924 38062
rect 35868 36484 35924 37996
rect 35868 36418 35924 36428
rect 35980 27636 36036 41916
rect 36204 40404 36260 40414
rect 36204 37044 36260 40348
rect 36204 36978 36260 36988
rect 35980 27570 36036 27580
rect 35756 24546 35812 24556
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 36316 21588 36372 47404
rect 36876 44996 36932 45006
rect 36764 43652 36820 43662
rect 36428 40964 36484 40974
rect 36428 21700 36484 40908
rect 36540 38612 36596 38622
rect 36540 38164 36596 38556
rect 36540 38098 36596 38108
rect 36764 38052 36820 43596
rect 36764 37986 36820 37996
rect 36540 37156 36596 37166
rect 36540 25172 36596 37100
rect 36876 28308 36932 44940
rect 40460 44436 40516 44446
rect 37436 43316 37492 43326
rect 37436 42644 37492 43260
rect 37436 42578 37492 42588
rect 40348 43316 40404 43326
rect 39452 42532 39508 42542
rect 39004 42084 39060 42094
rect 36876 28242 36932 28252
rect 36988 41972 37044 41982
rect 36988 27300 37044 41916
rect 37436 40964 37492 40974
rect 37100 40852 37156 40862
rect 37100 37828 37156 40796
rect 37100 37762 37156 37772
rect 37436 31108 37492 40908
rect 39004 40964 39060 42028
rect 38780 40404 38836 40414
rect 37436 31042 37492 31052
rect 38668 38836 38724 38846
rect 38668 32340 38724 38780
rect 36988 27234 37044 27244
rect 36540 25106 36596 25116
rect 36428 21634 36484 21644
rect 36316 21522 36372 21532
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 29372 11442 29428 11452
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 10220 35488 11732
rect 38668 11396 38724 32284
rect 38780 36708 38836 40348
rect 38780 16660 38836 36652
rect 39004 31780 39060 40908
rect 39004 31714 39060 31724
rect 38780 16594 38836 16604
rect 39452 16324 39508 42476
rect 39452 16258 39508 16268
rect 40348 13188 40404 43260
rect 40460 23268 40516 44380
rect 40460 23202 40516 23212
rect 40348 13122 40404 13132
rect 38668 11330 38724 11340
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 22848 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__155__I
timestamp 1663859327
transform 1 0 10976 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__A1
timestamp 1663859327
transform 1 0 15792 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__156__A2
timestamp 1663859327
transform -1 0 20384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__A1
timestamp 1663859327
transform -1 0 32816 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__157__A2
timestamp 1663859327
transform 1 0 32144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__I
timestamp 1663859327
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__A1
timestamp 1663859327
transform -1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__A2
timestamp 1663859327
transform -1 0 11312 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__A3
timestamp 1663859327
transform -1 0 12656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__A4
timestamp 1663859327
transform -1 0 11760 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__A1
timestamp 1663859327
transform 1 0 39088 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__A2
timestamp 1663859327
transform 1 0 37856 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__A3
timestamp 1663859327
transform 1 0 38640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__161__A4
timestamp 1663859327
transform 1 0 38192 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__A1
timestamp 1663859327
transform -1 0 7840 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__A3
timestamp 1663859327
transform -1 0 7392 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__A1
timestamp 1663859327
transform 1 0 28896 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__A2
timestamp 1663859327
transform 1 0 29904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__A3
timestamp 1663859327
transform -1 0 26656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__A4
timestamp 1663859327
transform 1 0 25088 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__A1
timestamp 1663859327
transform -1 0 23632 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__164__A2
timestamp 1663859327
transform -1 0 22624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__A1
timestamp 1663859327
transform 1 0 35728 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__A2
timestamp 1663859327
transform -1 0 35056 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__A3
timestamp 1663859327
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__165__A4
timestamp 1663859327
transform 1 0 35728 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__A1
timestamp 1663859327
transform 1 0 39088 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__A2
timestamp 1663859327
transform 1 0 38640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__A3
timestamp 1663859327
transform 1 0 38192 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__A4
timestamp 1663859327
transform 1 0 37408 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__I
timestamp 1663859327
transform 1 0 8960 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__A1
timestamp 1663859327
transform -1 0 20832 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__A2
timestamp 1663859327
transform -1 0 17920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__A3
timestamp 1663859327
transform -1 0 17808 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__A4
timestamp 1663859327
transform 1 0 17248 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A1
timestamp 1663859327
transform -1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A2
timestamp 1663859327
transform 1 0 13216 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A3
timestamp 1663859327
transform 1 0 13664 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A4
timestamp 1663859327
transform -1 0 17360 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__170__A1
timestamp 1663859327
transform -1 0 16240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__A1
timestamp 1663859327
transform 1 0 37744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__171__A4
timestamp 1663859327
transform 1 0 37408 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I
timestamp 1663859327
transform -1 0 3808 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__I
timestamp 1663859327
transform 1 0 7952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__A1
timestamp 1663859327
transform 1 0 35728 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__174__A2
timestamp 1663859327
transform 1 0 39536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__175__I
timestamp 1663859327
transform -1 0 2240 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__A1
timestamp 1663859327
transform 1 0 39200 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__176__A2
timestamp 1663859327
transform 1 0 39648 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__I
timestamp 1663859327
transform -1 0 13216 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__A1
timestamp 1663859327
transform -1 0 3136 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__178__A2
timestamp 1663859327
transform -1 0 2688 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__179__I
timestamp 1663859327
transform 1 0 16352 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__A1
timestamp 1663859327
transform 1 0 29680 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__A2
timestamp 1663859327
transform 1 0 30128 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__I
timestamp 1663859327
transform -1 0 10304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__I
timestamp 1663859327
transform -1 0 2464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__A1
timestamp 1663859327
transform 1 0 40096 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__183__A2
timestamp 1663859327
transform 1 0 40544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__A1
timestamp 1663859327
transform 1 0 32816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__A2
timestamp 1663859327
transform 1 0 32144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__I
timestamp 1663859327
transform -1 0 25760 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__A1
timestamp 1663859327
transform 1 0 33936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__187__A2
timestamp 1663859327
transform 1 0 34832 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__A1
timestamp 1663859327
transform -1 0 27104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__189__A2
timestamp 1663859327
transform -1 0 26656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__190__I
timestamp 1663859327
transform -1 0 6832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__A1
timestamp 1663859327
transform -1 0 2016 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__191__A2
timestamp 1663859327
transform -1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__I
timestamp 1663859327
transform -1 0 12656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__A1
timestamp 1663859327
transform -1 0 8288 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__A2
timestamp 1663859327
transform 1 0 7168 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__I
timestamp 1663859327
transform -1 0 11088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__A1
timestamp 1663859327
transform 1 0 37856 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__A2
timestamp 1663859327
transform 1 0 37520 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__I
timestamp 1663859327
transform -1 0 11760 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__A1
timestamp 1663859327
transform -1 0 12320 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__A2
timestamp 1663859327
transform -1 0 4704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A1
timestamp 1663859327
transform -1 0 6384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A2
timestamp 1663859327
transform 1 0 6608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__A4
timestamp 1663859327
transform -1 0 7728 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__A1
timestamp 1663859327
transform -1 0 15008 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__A2
timestamp 1663859327
transform -1 0 15680 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A1
timestamp 1663859327
transform -1 0 25760 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A2
timestamp 1663859327
transform -1 0 23520 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A3
timestamp 1663859327
transform -1 0 24976 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__A1
timestamp 1663859327
transform -1 0 23520 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__I
timestamp 1663859327
transform -1 0 6384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I0
timestamp 1663859327
transform 1 0 33936 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I1
timestamp 1663859327
transform 1 0 16688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I2
timestamp 1663859327
transform 1 0 35504 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I3
timestamp 1663859327
transform 1 0 5600 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__S0
timestamp 1663859327
transform 1 0 35952 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__S1
timestamp 1663859327
transform 1 0 36400 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__I
timestamp 1663859327
transform 1 0 9744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I0
timestamp 1663859327
transform 1 0 9744 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I1
timestamp 1663859327
transform -1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I2
timestamp 1663859327
transform 1 0 4032 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__I3
timestamp 1663859327
transform 1 0 4480 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__S0
timestamp 1663859327
transform -1 0 8736 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__S1
timestamp 1663859327
transform -1 0 9520 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I0
timestamp 1663859327
transform -1 0 7392 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I1
timestamp 1663859327
transform 1 0 8512 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I2
timestamp 1663859327
transform -1 0 9968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__I3
timestamp 1663859327
transform -1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__S0
timestamp 1663859327
transform -1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__S1
timestamp 1663859327
transform -1 0 7840 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__A1
timestamp 1663859327
transform 1 0 3584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__A2
timestamp 1663859327
transform -1 0 4256 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__I
timestamp 1663859327
transform 1 0 22400 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__I
timestamp 1663859327
transform 1 0 19712 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__A1
timestamp 1663859327
transform 1 0 39984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__A2
timestamp 1663859327
transform 1 0 39536 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__A1
timestamp 1663859327
transform -1 0 11312 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__A2
timestamp 1663859327
transform 1 0 15568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__A3
timestamp 1663859327
transform -1 0 14560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__I
timestamp 1663859327
transform -1 0 7840 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__I
timestamp 1663859327
transform 1 0 40880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__A1
timestamp 1663859327
transform 1 0 33488 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__A2
timestamp 1663859327
transform -1 0 34160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__A1
timestamp 1663859327
transform -1 0 5152 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__A2
timestamp 1663859327
transform 1 0 5824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__I
timestamp 1663859327
transform -1 0 31248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__A1
timestamp 1663859327
transform 1 0 38752 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__A2
timestamp 1663859327
transform 1 0 38304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__I
timestamp 1663859327
transform -1 0 2912 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__A1
timestamp 1663859327
transform -1 0 19264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__A2
timestamp 1663859327
transform -1 0 17136 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__A1
timestamp 1663859327
transform -1 0 3360 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__A2
timestamp 1663859327
transform 1 0 7056 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__A1
timestamp 1663859327
transform -1 0 4256 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__A2
timestamp 1663859327
transform -1 0 3808 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I
timestamp 1663859327
transform -1 0 5600 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__A1
timestamp 1663859327
transform -1 0 5152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__A2
timestamp 1663859327
transform -1 0 4256 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__A1
timestamp 1663859327
transform 1 0 32816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__A2
timestamp 1663859327
transform 1 0 33488 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__A3
timestamp 1663859327
transform 1 0 32368 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__B1
timestamp 1663859327
transform -1 0 32144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__B2
timestamp 1663859327
transform 1 0 35280 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__A1
timestamp 1663859327
transform -1 0 7168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__A2
timestamp 1663859327
transform -1 0 5376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__B
timestamp 1663859327
transform 1 0 6048 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__A1
timestamp 1663859327
transform -1 0 4704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__A2
timestamp 1663859327
transform -1 0 5600 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__A1
timestamp 1663859327
transform -1 0 23968 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__A2
timestamp 1663859327
transform 1 0 34832 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__I
timestamp 1663859327
transform -1 0 6048 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__I
timestamp 1663859327
transform -1 0 15456 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__A1
timestamp 1663859327
transform 1 0 10528 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__A2
timestamp 1663859327
transform 1 0 12544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__A1
timestamp 1663859327
transform 1 0 8848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__A2
timestamp 1663859327
transform 1 0 8400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I0
timestamp 1663859327
transform 1 0 37520 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__I1
timestamp 1663859327
transform 1 0 38416 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__S
timestamp 1663859327
transform 1 0 36624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__A1
timestamp 1663859327
transform -1 0 20160 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__A2
timestamp 1663859327
transform -1 0 18256 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__A3
timestamp 1663859327
transform -1 0 18816 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__A1
timestamp 1663859327
transform 1 0 40544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__A2
timestamp 1663859327
transform 1 0 40096 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__A1
timestamp 1663859327
transform 1 0 9296 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__A2
timestamp 1663859327
transform 1 0 8848 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__A3
timestamp 1663859327
transform 1 0 8064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__A1
timestamp 1663859327
transform -1 0 16128 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__A2
timestamp 1663859327
transform -1 0 14672 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__B
timestamp 1663859327
transform -1 0 18368 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__A2
timestamp 1663859327
transform 1 0 36400 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__A3
timestamp 1663859327
transform 1 0 36624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__B2
timestamp 1663859327
transform 1 0 35728 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__A1
timestamp 1663859327
transform -1 0 28000 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__A2
timestamp 1663859327
transform -1 0 28896 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__I
timestamp 1663859327
transform -1 0 21280 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__A1
timestamp 1663859327
transform 1 0 38864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__A2
timestamp 1663859327
transform 1 0 39200 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__B
timestamp 1663859327
transform 1 0 39648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__A1
timestamp 1663859327
transform -1 0 4704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__A2
timestamp 1663859327
transform -1 0 5936 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__I
timestamp 1663859327
transform -1 0 15232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__A1
timestamp 1663859327
transform 1 0 35280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__A2
timestamp 1663859327
transform -1 0 34608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A1
timestamp 1663859327
transform -1 0 19712 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A2
timestamp 1663859327
transform -1 0 19264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__A3
timestamp 1663859327
transform -1 0 21728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__A1
timestamp 1663859327
transform -1 0 4256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__248__A2
timestamp 1663859327
transform -1 0 3136 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__249__I
timestamp 1663859327
transform -1 0 7392 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__250__I
timestamp 1663859327
transform 1 0 13552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__251__I
timestamp 1663859327
transform 1 0 26880 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__A1
timestamp 1663859327
transform 1 0 35952 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__A2
timestamp 1663859327
transform 1 0 36176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__A1
timestamp 1663859327
transform 1 0 37072 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__A2
timestamp 1663859327
transform 1 0 37408 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__A1
timestamp 1663859327
transform -1 0 5152 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__A2
timestamp 1663859327
transform -1 0 6048 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__A1
timestamp 1663859327
transform -1 0 24752 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__A2
timestamp 1663859327
transform -1 0 24416 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__A3
timestamp 1663859327
transform 1 0 20832 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__I
timestamp 1663859327
transform 1 0 31920 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__A1
timestamp 1663859327
transform 1 0 25984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__A2
timestamp 1663859327
transform -1 0 25312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__A1
timestamp 1663859327
transform 1 0 30688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__A2
timestamp 1663859327
transform -1 0 33712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__A3
timestamp 1663859327
transform 1 0 33488 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I
timestamp 1663859327
transform 1 0 28448 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__A1
timestamp 1663859327
transform 1 0 37296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__A2
timestamp 1663859327
transform 1 0 33040 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__A3
timestamp 1663859327
transform 1 0 34832 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__B
timestamp 1663859327
transform 1 0 34384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__A1
timestamp 1663859327
transform 1 0 38864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__A2
timestamp 1663859327
transform 1 0 35728 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__A3
timestamp 1663859327
transform 1 0 34832 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__A1
timestamp 1663859327
transform 1 0 31696 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__A2
timestamp 1663859327
transform 1 0 33040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__B
timestamp 1663859327
transform -1 0 31472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__A1
timestamp 1663859327
transform 1 0 10640 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__A2
timestamp 1663859327
transform -1 0 10864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__A3
timestamp 1663859327
transform 1 0 10192 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__A1
timestamp 1663859327
transform -1 0 23072 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__A2
timestamp 1663859327
transform 1 0 21952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__A1
timestamp 1663859327
transform -1 0 16240 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__A2
timestamp 1663859327
transform -1 0 9968 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__B
timestamp 1663859327
transform -1 0 11648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__I
timestamp 1663859327
transform -1 0 14896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__A1
timestamp 1663859327
transform -1 0 13664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__A3
timestamp 1663859327
transform 1 0 10640 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__A1
timestamp 1663859327
transform -1 0 19152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__A2
timestamp 1663859327
transform 1 0 18480 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__A1
timestamp 1663859327
transform 1 0 41440 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__A2
timestamp 1663859327
transform 1 0 40432 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__A2
timestamp 1663859327
transform 1 0 40208 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__270__B2
timestamp 1663859327
transform 1 0 38416 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__A1
timestamp 1663859327
transform 1 0 37968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__A2
timestamp 1663859327
transform -1 0 8288 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__271__B
timestamp 1663859327
transform -1 0 9072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__A1
timestamp 1663859327
transform -1 0 27552 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__272__A2
timestamp 1663859327
transform -1 0 28448 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__A1
timestamp 1663859327
transform 1 0 34384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__274__A2
timestamp 1663859327
transform 1 0 33488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__A1
timestamp 1663859327
transform -1 0 25760 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__A2
timestamp 1663859327
transform -1 0 27552 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__B1
timestamp 1663859327
transform -1 0 24864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__275__B2
timestamp 1663859327
transform 1 0 29344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__A1
timestamp 1663859327
transform -1 0 32816 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__A2
timestamp 1663859327
transform -1 0 32816 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__B1
timestamp 1663859327
transform 1 0 36848 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__B2
timestamp 1663859327
transform 1 0 37296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__276__C
timestamp 1663859327
transform 1 0 36400 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__277__A1
timestamp 1663859327
transform 1 0 40208 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__277__A2
timestamp 1663859327
transform 1 0 40656 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__A1
timestamp 1663859327
transform 1 0 32368 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__278__A2
timestamp 1663859327
transform 1 0 29456 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__A1
timestamp 1663859327
transform -1 0 2688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__A2
timestamp 1663859327
transform -1 0 3808 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__279__B
timestamp 1663859327
transform -1 0 2240 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__A1
timestamp 1663859327
transform -1 0 6944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__280__A2
timestamp 1663859327
transform -1 0 7840 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__A1
timestamp 1663859327
transform -1 0 17024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__A2
timestamp 1663859327
transform 1 0 17696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__A3
timestamp 1663859327
transform 1 0 16128 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__281__B
timestamp 1663859327
transform 1 0 15680 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__A1
timestamp 1663859327
transform -1 0 14112 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__A2
timestamp 1663859327
transform -1 0 12096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__282__B
timestamp 1663859327
transform -1 0 10416 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__283__A1
timestamp 1663859327
transform -1 0 3584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__283__A2
timestamp 1663859327
transform -1 0 4032 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A1
timestamp 1663859327
transform 1 0 32144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__A2
timestamp 1663859327
transform -1 0 32816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__B1
timestamp 1663859327
transform 1 0 30352 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__B2
timestamp 1663859327
transform 1 0 30800 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__284__C
timestamp 1663859327
transform 1 0 31696 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__A1
timestamp 1663859327
transform -1 0 3360 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__285__A2
timestamp 1663859327
transform -1 0 2912 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__A1
timestamp 1663859327
transform 1 0 31136 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__A2
timestamp 1663859327
transform 1 0 35728 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__286__B
timestamp 1663859327
transform 1 0 35280 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A1
timestamp 1663859327
transform 1 0 35280 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__A2
timestamp 1663859327
transform 1 0 34384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__287__B
timestamp 1663859327
transform 1 0 36176 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__I0
timestamp 1663859327
transform -1 0 7392 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__I1
timestamp 1663859327
transform -1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__289__S
timestamp 1663859327
transform -1 0 8176 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A1
timestamp 1663859327
transform 1 0 39312 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A2
timestamp 1663859327
transform 1 0 40656 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__290__A3
timestamp 1663859327
transform 1 0 39760 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__291__A2
timestamp 1663859327
transform 1 0 38752 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__292__I
timestamp 1663859327
transform 1 0 34832 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A1
timestamp 1663859327
transform -1 0 14336 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__293__A2
timestamp 1663859327
transform -1 0 14784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__A1
timestamp 1663859327
transform 1 0 37408 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__294__A2
timestamp 1663859327
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__A1
timestamp 1663859327
transform 1 0 39312 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__A2
timestamp 1663859327
transform 1 0 36176 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__295__C
timestamp 1663859327
transform -1 0 37184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A1
timestamp 1663859327
transform -1 0 2912 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__A2
timestamp 1663859327
transform -1 0 3808 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__296__B
timestamp 1663859327
transform -1 0 4256 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A1
timestamp 1663859327
transform 1 0 31696 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__A2
timestamp 1663859327
transform 1 0 34384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__297__B
timestamp 1663859327
transform 1 0 33936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__A1
timestamp 1663859327
transform -1 0 4928 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__A2
timestamp 1663859327
transform 1 0 6720 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__B1
timestamp 1663859327
transform -1 0 4480 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__B2
timestamp 1663859327
transform -1 0 5152 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__C1
timestamp 1663859327
transform -1 0 5824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__298__C2
timestamp 1663859327
transform 1 0 5152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__A1
timestamp 1663859327
transform -1 0 9856 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__299__A2
timestamp 1663859327
transform -1 0 7840 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__A1
timestamp 1663859327
transform -1 0 29680 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__B1
timestamp 1663859327
transform 1 0 30576 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__B2
timestamp 1663859327
transform -1 0 27104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__300__C
timestamp 1663859327
transform 1 0 31472 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__A1
timestamp 1663859327
transform 1 0 37072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__A2
timestamp 1663859327
transform 1 0 36624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__A3
timestamp 1663859327
transform 1 0 36176 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__301__A4
timestamp 1663859327
transform 1 0 34384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A1
timestamp 1663859327
transform 1 0 38864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A2
timestamp 1663859327
transform -1 0 9856 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A3
timestamp 1663859327
transform -1 0 10752 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__302__A4
timestamp 1663859327
transform 1 0 37968 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__A1
timestamp 1663859327
transform -1 0 5152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__303__A2
timestamp 1663859327
transform -1 0 4704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A1
timestamp 1663859327
transform 1 0 29792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A2
timestamp 1663859327
transform -1 0 22624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A3
timestamp 1663859327
transform -1 0 31024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__304__A4
timestamp 1663859327
transform -1 0 28000 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A1
timestamp 1663859327
transform -1 0 5936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__A2
timestamp 1663859327
transform -1 0 4704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__305__B
timestamp 1663859327
transform -1 0 5600 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__A1
timestamp 1663859327
transform 1 0 35280 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__A2
timestamp 1663859327
transform 1 0 34384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__B1
timestamp 1663859327
transform 1 0 33936 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__B2
timestamp 1663859327
transform 1 0 34832 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__306__C
timestamp 1663859327
transform 1 0 33488 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__A1
timestamp 1663859327
transform 1 0 39760 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__A2
timestamp 1663859327
transform 1 0 39312 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__308__B
timestamp 1663859327
transform 1 0 38304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__A1
timestamp 1663859327
transform 1 0 31472 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__A2
timestamp 1663859327
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__309__B
timestamp 1663859327
transform 1 0 33488 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__A1
timestamp 1663859327
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__310__B1
timestamp 1663859327
transform -1 0 9968 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__A1
timestamp 1663859327
transform 1 0 39648 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__A2
timestamp 1663859327
transform 1 0 39200 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__B
timestamp 1663859327
transform 1 0 38304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__311__C
timestamp 1663859327
transform 1 0 38752 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A1
timestamp 1663859327
transform 1 0 3136 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__312__A2
timestamp 1663859327
transform -1 0 4704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__313__I
timestamp 1663859327
transform -1 0 24080 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__314__I
timestamp 1663859327
transform 1 0 6272 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__A1
timestamp 1663859327
transform 1 0 38752 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__A2
timestamp 1663859327
transform -1 0 38528 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__B
timestamp 1663859327
transform 1 0 37520 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__315__C
timestamp 1663859327
transform -1 0 38080 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A1
timestamp 1663859327
transform -1 0 30464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__316__A2
timestamp 1663859327
transform -1 0 31472 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__318__I
timestamp 1663859327
transform -1 0 30576 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__A1
timestamp 1663859327
transform -1 0 2464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__A2
timestamp 1663859327
transform -1 0 3584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__B
timestamp 1663859327
transform -1 0 4032 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__319__C
timestamp 1663859327
transform -1 0 2912 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__A1
timestamp 1663859327
transform 1 0 37072 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__320__A2
timestamp 1663859327
transform 1 0 38416 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__321__I
timestamp 1663859327
transform 1 0 28000 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__A1
timestamp 1663859327
transform -1 0 26208 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__A2
timestamp 1663859327
transform -1 0 23968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__B
timestamp 1663859327
transform -1 0 22064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__322__C
timestamp 1663859327
transform -1 0 24528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__323__A1
timestamp 1663859327
transform -1 0 15568 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__324__I
timestamp 1663859327
transform -1 0 8736 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__CLK
timestamp 1663859327
transform 1 0 35504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__325__D
timestamp 1663859327
transform 1 0 35056 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__CLK
timestamp 1663859327
transform 1 0 8064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__326__D
timestamp 1663859327
transform -1 0 28448 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__CLK
timestamp 1663859327
transform 1 0 6720 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__327__D
timestamp 1663859327
transform -1 0 7840 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__CLK
timestamp 1663859327
transform 1 0 6496 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__328__D
timestamp 1663859327
transform -1 0 6272 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__CLK
timestamp 1663859327
transform 1 0 6272 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__329__D
timestamp 1663859327
transform -1 0 5936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__CLK
timestamp 1663859327
transform 1 0 5600 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__330__D
timestamp 1663859327
transform -1 0 7280 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__CLK
timestamp 1663859327
transform 1 0 8512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__331__D
timestamp 1663859327
transform -1 0 10304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__332__CLK
timestamp 1663859327
transform 1 0 5824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__CLK
timestamp 1663859327
transform 1 0 6272 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__333__D
timestamp 1663859327
transform -1 0 7728 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__334__CLK
timestamp 1663859327
transform 1 0 7392 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__CLK
timestamp 1663859327
transform 1 0 8400 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__335__D
timestamp 1663859327
transform -1 0 10080 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__CLK
timestamp 1663859327
transform 1 0 9744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__336__D
timestamp 1663859327
transform -1 0 23072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__CLK
timestamp 1663859327
transform -1 0 14224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__337__D
timestamp 1663859327
transform -1 0 17920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__CLK
timestamp 1663859327
transform 1 0 6160 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__338__D
timestamp 1663859327
transform -1 0 7280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__CLK
timestamp 1663859327
transform 1 0 33936 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__339__D
timestamp 1663859327
transform -1 0 33712 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__CLK
timestamp 1663859327
transform 1 0 6272 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__340__D
timestamp 1663859327
transform -1 0 6832 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__CLK
timestamp 1663859327
transform 1 0 11536 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__341__D
timestamp 1663859327
transform -1 0 12544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__CLK
timestamp 1663859327
transform 1 0 6720 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__342__D
timestamp 1663859327
transform -1 0 9072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__CLK
timestamp 1663859327
transform 1 0 35952 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__343__D
timestamp 1663859327
transform 1 0 35504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__344__CLK
timestamp 1663859327
transform 1 0 7952 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__CLK
timestamp 1663859327
transform 1 0 10192 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__345__D
timestamp 1663859327
transform -1 0 11312 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__CLK
timestamp 1663859327
transform 1 0 6160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__346__D
timestamp 1663859327
transform -1 0 8288 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__CLK
timestamp 1663859327
transform 1 0 17584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__347__D
timestamp 1663859327
transform 1 0 32816 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__CLK
timestamp 1663859327
transform 1 0 11984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__348__D
timestamp 1663859327
transform -1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__CLK
timestamp 1663859327
transform 1 0 7504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__349__D
timestamp 1663859327
transform -1 0 6496 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__CLK
timestamp 1663859327
transform 1 0 6720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__350__D
timestamp 1663859327
transform -1 0 7280 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__351__CLK
timestamp 1663859327
transform 1 0 4928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__CLK
timestamp 1663859327
transform 1 0 4480 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__352__D
timestamp 1663859327
transform -1 0 5600 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__CLK
timestamp 1663859327
transform 1 0 14112 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__353__D
timestamp 1663859327
transform -1 0 15120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__CLK
timestamp 1663859327
transform 1 0 9296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__354__D
timestamp 1663859327
transform -1 0 12208 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__CLK
timestamp 1663859327
transform 1 0 8960 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__355__D
timestamp 1663859327
transform -1 0 8736 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__CLK
timestamp 1663859327
transform 1 0 34384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__356__D
timestamp 1663859327
transform 1 0 35280 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__CLK
timestamp 1663859327
transform -1 0 5152 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__357__D
timestamp 1663859327
transform -1 0 6048 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__CLK
timestamp 1663859327
transform 1 0 34832 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__358__D
timestamp 1663859327
transform 1 0 35728 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__359__CLK
timestamp 1663859327
transform 1 0 36848 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__CLK
timestamp 1663859327
transform 1 0 37856 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__360__D
timestamp 1663859327
transform 1 0 35280 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__CLK
timestamp 1663859327
transform 1 0 33936 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__361__D
timestamp 1663859327
transform 1 0 36176 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__CLK
timestamp 1663859327
transform 1 0 33040 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__362__D
timestamp 1663859327
transform 1 0 28672 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__CLK
timestamp 1663859327
transform 1 0 4704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__363__D
timestamp 1663859327
transform -1 0 4480 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__CLK
timestamp 1663859327
transform 1 0 6608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__364__D
timestamp 1663859327
transform -1 0 4256 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__CLK
timestamp 1663859327
transform -1 0 3808 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__365__D
timestamp 1663859327
transform -1 0 3360 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__CLK
timestamp 1663859327
transform 1 0 6048 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__366__D
timestamp 1663859327
transform 1 0 37744 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__CLK
timestamp 1663859327
transform 1 0 11984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__367__D
timestamp 1663859327
transform -1 0 12992 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__CLK
timestamp 1663859327
transform 1 0 8176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__368__D
timestamp 1663859327
transform -1 0 9856 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__CLK
timestamp 1663859327
transform 1 0 8400 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__369__D
timestamp 1663859327
transform 1 0 36176 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__CLK
timestamp 1663859327
transform 1 0 9296 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__370__D
timestamp 1663859327
transform 1 0 32592 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__440__I
timestamp 1663859327
transform 1 0 3808 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__441__I
timestamp 1663859327
transform 1 0 9520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1663859327
transform -1 0 2016 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1663859327
transform -1 0 47600 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1663859327
transform -1 0 47376 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1663859327
transform -1 0 36512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1663859327
transform -1 0 11984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1663859327
transform -1 0 1904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1663859327
transform -1 0 18704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1663859327
transform 1 0 41328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output9_I
timestamp 1663859327
transform 1 0 4032 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output10_I
timestamp 1663859327
transform -1 0 7392 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output11_I
timestamp 1663859327
transform 1 0 41776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output12_I
timestamp 1663859327
transform -1 0 2464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output13_I
timestamp 1663859327
transform 1 0 3472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output14_I
timestamp 1663859327
transform -1 0 4368 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output15_I
timestamp 1663859327
transform 1 0 40096 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1568 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 3248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23
timestamp 1663859327
transform 1 0 3920 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 4368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37
timestamp 1663859327
transform 1 0 5488 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 6048 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58
timestamp 1663859327
transform 1 0 7840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_66 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 8736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_72
timestamp 1663859327
transform 1 0 9408 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_77
timestamp 1663859327
transform 1 0 9968 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_95
timestamp 1663859327
transform 1 0 11984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_103
timestamp 1663859327
transform 1 0 12880 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_107
timestamp 1663859327
transform 1 0 13328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_119
timestamp 1663859327
transform 1 0 14672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_131
timestamp 1663859327
transform 1 0 16016 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_139
timestamp 1663859327
transform 1 0 16912 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_142
timestamp 1663859327
transform 1 0 17248 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_144
timestamp 1663859327
transform 1 0 17472 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_149
timestamp 1663859327
transform 1 0 18032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_155
timestamp 1663859327
transform 1 0 18704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_163
timestamp 1663859327
transform 1 0 19600 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_171
timestamp 1663859327
transform 1 0 20496 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_177
timestamp 1663859327
transform 1 0 21168 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_182
timestamp 1663859327
transform 1 0 21728 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_190
timestamp 1663859327
transform 1 0 22624 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_192
timestamp 1663859327
transform 1 0 22848 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_197
timestamp 1663859327
transform 1 0 23408 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_205
timestamp 1663859327
transform 1 0 24304 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_209
timestamp 1663859327
transform 1 0 24752 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_212
timestamp 1663859327
transform 1 0 25088 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_220
timestamp 1663859327
transform 1 0 25984 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_222
timestamp 1663859327
transform 1 0 26208 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_227
timestamp 1663859327
transform 1 0 26768 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_243
timestamp 1663859327
transform 1 0 28560 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_247
timestamp 1663859327
transform 1 0 29008 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_252
timestamp 1663859327
transform 1 0 29568 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_268
timestamp 1663859327
transform 1 0 31360 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_270
timestamp 1663859327
transform 1 0 31584 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_275
timestamp 1663859327
transform 1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_279
timestamp 1663859327
transform 1 0 32592 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_282
timestamp 1663859327
transform 1 0 32928 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_298
timestamp 1663859327
transform 1 0 34720 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_300
timestamp 1663859327
transform 1 0 34944 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_305
timestamp 1663859327
transform 1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_309
timestamp 1663859327
transform 1 0 35952 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_311
timestamp 1663859327
transform 1 0 36176 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_314
timestamp 1663859327
transform 1 0 36512 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_317
timestamp 1663859327
transform 1 0 36848 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_325
timestamp 1663859327
transform 1 0 37744 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_329
timestamp 1663859327
transform 1 0 38192 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_335
timestamp 1663859327
transform 1 0 38864 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_343
timestamp 1663859327
transform 1 0 39760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_347
timestamp 1663859327
transform 1 0 40208 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_349
timestamp 1663859327
transform 1 0 40432 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_352
timestamp 1663859327
transform 1 0 40768 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_357
timestamp 1663859327
transform 1 0 41328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_365
timestamp 1663859327
transform 1 0 42224 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_371
timestamp 1663859327
transform 1 0 42896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_383
timestamp 1663859327
transform 1 0 44240 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_387
timestamp 1663859327
transform 1 0 44688 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_395
timestamp 1663859327
transform 1 0 45584 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_401
timestamp 1663859327
transform 1 0 46256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_405
timestamp 1663859327
transform 1 0 46704 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_411
timestamp 1663859327
transform 1 0 47376 0 1 3136
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_419
timestamp 1663859327
transform 1 0 48272 0 1 3136
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_2
timestamp 1663859327
transform 1 0 1568 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_7
timestamp 1663859327
transform 1 0 2128 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_13 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 2800 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_45
timestamp 1663859327
transform 1 0 6384 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_1_61
timestamp 1663859327
transform 1 0 8176 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_69
timestamp 1663859327
transform 1 0 9072 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_73 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 9520 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_137
timestamp 1663859327
transform 1 0 16688 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_141
timestamp 1663859327
transform 1 0 17136 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_144
timestamp 1663859327
transform 1 0 17472 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_208
timestamp 1663859327
transform 1 0 24640 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_212
timestamp 1663859327
transform 1 0 25088 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_215
timestamp 1663859327
transform 1 0 25424 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_279
timestamp 1663859327
transform 1 0 32592 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_283
timestamp 1663859327
transform 1 0 33040 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_1_286
timestamp 1663859327
transform 1 0 33376 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_350
timestamp 1663859327
transform 1 0 40544 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_354
timestamp 1663859327
transform 1 0 40992 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_1_357
timestamp 1663859327
transform 1 0 41328 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_1_389
timestamp 1663859327
transform 1 0 44912 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_1_405
timestamp 1663859327
transform 1 0 46704 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_409
timestamp 1663859327
transform 1 0 47152 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_1_413
timestamp 1663859327
transform 1 0 47600 0 -1 4704
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_1_419
timestamp 1663859327
transform 1 0 48272 0 -1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_2_2
timestamp 1663859327
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_34
timestamp 1663859327
transform 1 0 5152 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_37
timestamp 1663859327
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_101
timestamp 1663859327
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_105
timestamp 1663859327
transform 1 0 13104 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_108
timestamp 1663859327
transform 1 0 13440 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_172
timestamp 1663859327
transform 1 0 20608 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_176
timestamp 1663859327
transform 1 0 21056 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_179
timestamp 1663859327
transform 1 0 21392 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_243
timestamp 1663859327
transform 1 0 28560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_247
timestamp 1663859327
transform 1 0 29008 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_250
timestamp 1663859327
transform 1 0 29344 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_314
timestamp 1663859327
transform 1 0 36512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_318
timestamp 1663859327
transform 1 0 36960 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_2_321
timestamp 1663859327
transform 1 0 37296 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_385
timestamp 1663859327
transform 1 0 44464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_2_389
timestamp 1663859327
transform 1 0 44912 0 1 4704
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_2_392
timestamp 1663859327
transform 1 0 45248 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_2_408
timestamp 1663859327
transform 1 0 47040 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_2_416
timestamp 1663859327
transform 1 0 47936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_2
timestamp 1663859327
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_66
timestamp 1663859327
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_70
timestamp 1663859327
transform 1 0 9184 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_73
timestamp 1663859327
transform 1 0 9520 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_137
timestamp 1663859327
transform 1 0 16688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_141
timestamp 1663859327
transform 1 0 17136 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_144
timestamp 1663859327
transform 1 0 17472 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_208
timestamp 1663859327
transform 1 0 24640 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_212
timestamp 1663859327
transform 1 0 25088 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_215
timestamp 1663859327
transform 1 0 25424 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_279
timestamp 1663859327
transform 1 0 32592 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_283
timestamp 1663859327
transform 1 0 33040 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_3_286
timestamp 1663859327
transform 1 0 33376 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_350
timestamp 1663859327
transform 1 0 40544 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_354
timestamp 1663859327
transform 1 0 40992 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_3_357
timestamp 1663859327
transform 1 0 41328 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_3_389
timestamp 1663859327
transform 1 0 44912 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_3_405
timestamp 1663859327
transform 1 0 46704 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_3_413
timestamp 1663859327
transform 1 0 47600 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_3_417
timestamp 1663859327
transform 1 0 48048 0 -1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_3_419
timestamp 1663859327
transform 1 0 48272 0 -1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_4_2
timestamp 1663859327
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_34
timestamp 1663859327
transform 1 0 5152 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_37
timestamp 1663859327
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_101
timestamp 1663859327
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_105
timestamp 1663859327
transform 1 0 13104 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_108
timestamp 1663859327
transform 1 0 13440 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_172
timestamp 1663859327
transform 1 0 20608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_176
timestamp 1663859327
transform 1 0 21056 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_179
timestamp 1663859327
transform 1 0 21392 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_243
timestamp 1663859327
transform 1 0 28560 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_247
timestamp 1663859327
transform 1 0 29008 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_250
timestamp 1663859327
transform 1 0 29344 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_314
timestamp 1663859327
transform 1 0 36512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_318
timestamp 1663859327
transform 1 0 36960 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_4_321
timestamp 1663859327
transform 1 0 37296 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_385
timestamp 1663859327
transform 1 0 44464 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_389
timestamp 1663859327
transform 1 0 44912 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_4_392
timestamp 1663859327
transform 1 0 45248 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_4_408
timestamp 1663859327
transform 1 0 47040 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_4_412
timestamp 1663859327
transform 1 0 47488 0 1 6272
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_414
timestamp 1663859327
transform 1 0 47712 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_4_419
timestamp 1663859327
transform 1 0 48272 0 1 6272
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_2
timestamp 1663859327
transform 1 0 1568 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_7
timestamp 1663859327
transform 1 0 2128 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_73
timestamp 1663859327
transform 1 0 9520 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_137
timestamp 1663859327
transform 1 0 16688 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_141
timestamp 1663859327
transform 1 0 17136 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_144
timestamp 1663859327
transform 1 0 17472 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_208
timestamp 1663859327
transform 1 0 24640 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_212
timestamp 1663859327
transform 1 0 25088 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_215
timestamp 1663859327
transform 1 0 25424 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_279
timestamp 1663859327
transform 1 0 32592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_283
timestamp 1663859327
transform 1 0 33040 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_5_286
timestamp 1663859327
transform 1 0 33376 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_350
timestamp 1663859327
transform 1 0 40544 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_354
timestamp 1663859327
transform 1 0 40992 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_5_357
timestamp 1663859327
transform 1 0 41328 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_5_389
timestamp 1663859327
transform 1 0 44912 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_5_405
timestamp 1663859327
transform 1 0 46704 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_5_413
timestamp 1663859327
transform 1 0 47600 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_5_417
timestamp 1663859327
transform 1 0 48048 0 -1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_5_419
timestamp 1663859327
transform 1 0 48272 0 -1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_6_2
timestamp 1663859327
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_34
timestamp 1663859327
transform 1 0 5152 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_37
timestamp 1663859327
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_101
timestamp 1663859327
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_105
timestamp 1663859327
transform 1 0 13104 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_108
timestamp 1663859327
transform 1 0 13440 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_172
timestamp 1663859327
transform 1 0 20608 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_176
timestamp 1663859327
transform 1 0 21056 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_179
timestamp 1663859327
transform 1 0 21392 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_243
timestamp 1663859327
transform 1 0 28560 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_247
timestamp 1663859327
transform 1 0 29008 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_250
timestamp 1663859327
transform 1 0 29344 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_314
timestamp 1663859327
transform 1 0 36512 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_318
timestamp 1663859327
transform 1 0 36960 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_6_321
timestamp 1663859327
transform 1 0 37296 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_385
timestamp 1663859327
transform 1 0 44464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_389
timestamp 1663859327
transform 1 0 44912 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_6_392
timestamp 1663859327
transform 1 0 45248 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_6_408
timestamp 1663859327
transform 1 0 47040 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_6_412
timestamp 1663859327
transform 1 0 47488 0 1 7840
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_414
timestamp 1663859327
transform 1 0 47712 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_6_419
timestamp 1663859327
transform 1 0 48272 0 1 7840
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_2
timestamp 1663859327
transform 1 0 1568 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_7
timestamp 1663859327
transform 1 0 2128 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_73
timestamp 1663859327
transform 1 0 9520 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_137
timestamp 1663859327
transform 1 0 16688 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_141
timestamp 1663859327
transform 1 0 17136 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_144
timestamp 1663859327
transform 1 0 17472 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_208
timestamp 1663859327
transform 1 0 24640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_212
timestamp 1663859327
transform 1 0 25088 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_215
timestamp 1663859327
transform 1 0 25424 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_279
timestamp 1663859327
transform 1 0 32592 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_283
timestamp 1663859327
transform 1 0 33040 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_7_286
timestamp 1663859327
transform 1 0 33376 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_350
timestamp 1663859327
transform 1 0 40544 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_354
timestamp 1663859327
transform 1 0 40992 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_7_357
timestamp 1663859327
transform 1 0 41328 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_7_389
timestamp 1663859327
transform 1 0 44912 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_7_405
timestamp 1663859327
transform 1 0 46704 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_7_413
timestamp 1663859327
transform 1 0 47600 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_7_417
timestamp 1663859327
transform 1 0 48048 0 -1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_7_419
timestamp 1663859327
transform 1 0 48272 0 -1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_8_2
timestamp 1663859327
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_34
timestamp 1663859327
transform 1 0 5152 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_37
timestamp 1663859327
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_53
timestamp 1663859327
transform 1 0 7280 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_61
timestamp 1663859327
transform 1 0 8176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_71
timestamp 1663859327
transform 1 0 9296 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_75
timestamp 1663859327
transform 1 0 9744 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_8_91
timestamp 1663859327
transform 1 0 11536 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_99
timestamp 1663859327
transform 1 0 12432 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_103
timestamp 1663859327
transform 1 0 12880 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_105
timestamp 1663859327
transform 1 0 13104 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_108
timestamp 1663859327
transform 1 0 13440 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_172
timestamp 1663859327
transform 1 0 20608 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_176
timestamp 1663859327
transform 1 0 21056 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_179
timestamp 1663859327
transform 1 0 21392 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_243
timestamp 1663859327
transform 1 0 28560 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_247
timestamp 1663859327
transform 1 0 29008 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_250
timestamp 1663859327
transform 1 0 29344 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_314
timestamp 1663859327
transform 1 0 36512 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_318
timestamp 1663859327
transform 1 0 36960 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_8_321
timestamp 1663859327
transform 1 0 37296 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_385
timestamp 1663859327
transform 1 0 44464 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_389
timestamp 1663859327
transform 1 0 44912 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_8_392
timestamp 1663859327
transform 1 0 45248 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_8_408
timestamp 1663859327
transform 1 0 47040 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_8_412
timestamp 1663859327
transform 1 0 47488 0 1 9408
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_414
timestamp 1663859327
transform 1 0 47712 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_8_419
timestamp 1663859327
transform 1 0 48272 0 1 9408
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_2
timestamp 1663859327
transform 1 0 1568 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_7
timestamp 1663859327
transform 1 0 2128 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_73
timestamp 1663859327
transform 1 0 9520 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_137
timestamp 1663859327
transform 1 0 16688 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_141
timestamp 1663859327
transform 1 0 17136 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_144
timestamp 1663859327
transform 1 0 17472 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_208
timestamp 1663859327
transform 1 0 24640 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_212
timestamp 1663859327
transform 1 0 25088 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_215
timestamp 1663859327
transform 1 0 25424 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_279
timestamp 1663859327
transform 1 0 32592 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_283
timestamp 1663859327
transform 1 0 33040 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_9_286
timestamp 1663859327
transform 1 0 33376 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_350
timestamp 1663859327
transform 1 0 40544 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_354
timestamp 1663859327
transform 1 0 40992 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_9_357
timestamp 1663859327
transform 1 0 41328 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_9_389
timestamp 1663859327
transform 1 0 44912 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_9_405
timestamp 1663859327
transform 1 0 46704 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_9_413
timestamp 1663859327
transform 1 0 47600 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_9_417
timestamp 1663859327
transform 1 0 48048 0 -1 10976
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_9_419
timestamp 1663859327
transform 1 0 48272 0 -1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_10_2
timestamp 1663859327
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_34
timestamp 1663859327
transform 1 0 5152 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_37
timestamp 1663859327
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_101
timestamp 1663859327
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_105
timestamp 1663859327
transform 1 0 13104 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_108
timestamp 1663859327
transform 1 0 13440 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_172
timestamp 1663859327
transform 1 0 20608 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_176
timestamp 1663859327
transform 1 0 21056 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_179
timestamp 1663859327
transform 1 0 21392 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_243
timestamp 1663859327
transform 1 0 28560 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_247
timestamp 1663859327
transform 1 0 29008 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_250
timestamp 1663859327
transform 1 0 29344 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_314
timestamp 1663859327
transform 1 0 36512 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_318
timestamp 1663859327
transform 1 0 36960 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_10_321
timestamp 1663859327
transform 1 0 37296 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_385
timestamp 1663859327
transform 1 0 44464 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_10_389
timestamp 1663859327
transform 1 0 44912 0 1 10976
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_10_392
timestamp 1663859327
transform 1 0 45248 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_10_408
timestamp 1663859327
transform 1 0 47040 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_10_416
timestamp 1663859327
transform 1 0 47936 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_2
timestamp 1663859327
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_66
timestamp 1663859327
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_70
timestamp 1663859327
transform 1 0 9184 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_73
timestamp 1663859327
transform 1 0 9520 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_137
timestamp 1663859327
transform 1 0 16688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_141
timestamp 1663859327
transform 1 0 17136 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_144
timestamp 1663859327
transform 1 0 17472 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_208
timestamp 1663859327
transform 1 0 24640 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_212
timestamp 1663859327
transform 1 0 25088 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_215
timestamp 1663859327
transform 1 0 25424 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_279
timestamp 1663859327
transform 1 0 32592 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_283
timestamp 1663859327
transform 1 0 33040 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_11_286
timestamp 1663859327
transform 1 0 33376 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_11_350
timestamp 1663859327
transform 1 0 40544 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_354
timestamp 1663859327
transform 1 0 40992 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_11_357
timestamp 1663859327
transform 1 0 41328 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_11_389
timestamp 1663859327
transform 1 0 44912 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_11_405
timestamp 1663859327
transform 1 0 46704 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_11_413
timestamp 1663859327
transform 1 0 47600 0 -1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_11_419
timestamp 1663859327
transform 1 0 48272 0 -1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_12_2
timestamp 1663859327
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_34
timestamp 1663859327
transform 1 0 5152 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_37
timestamp 1663859327
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_101
timestamp 1663859327
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_105
timestamp 1663859327
transform 1 0 13104 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_108
timestamp 1663859327
transform 1 0 13440 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_172
timestamp 1663859327
transform 1 0 20608 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_176
timestamp 1663859327
transform 1 0 21056 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_179
timestamp 1663859327
transform 1 0 21392 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_243
timestamp 1663859327
transform 1 0 28560 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_247
timestamp 1663859327
transform 1 0 29008 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_250
timestamp 1663859327
transform 1 0 29344 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_314
timestamp 1663859327
transform 1 0 36512 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_318
timestamp 1663859327
transform 1 0 36960 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_12_321
timestamp 1663859327
transform 1 0 37296 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_385
timestamp 1663859327
transform 1 0 44464 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_389
timestamp 1663859327
transform 1 0 44912 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_12_392
timestamp 1663859327
transform 1 0 45248 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_12_408
timestamp 1663859327
transform 1 0 47040 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_12_412
timestamp 1663859327
transform 1 0 47488 0 1 12544
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_414
timestamp 1663859327
transform 1 0 47712 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_12_419
timestamp 1663859327
transform 1 0 48272 0 1 12544
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_2
timestamp 1663859327
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_66
timestamp 1663859327
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_70
timestamp 1663859327
transform 1 0 9184 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_73
timestamp 1663859327
transform 1 0 9520 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_137
timestamp 1663859327
transform 1 0 16688 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_141
timestamp 1663859327
transform 1 0 17136 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_144
timestamp 1663859327
transform 1 0 17472 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_208
timestamp 1663859327
transform 1 0 24640 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_212
timestamp 1663859327
transform 1 0 25088 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_215
timestamp 1663859327
transform 1 0 25424 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_279
timestamp 1663859327
transform 1 0 32592 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_283
timestamp 1663859327
transform 1 0 33040 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_13_286
timestamp 1663859327
transform 1 0 33376 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_350
timestamp 1663859327
transform 1 0 40544 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_354
timestamp 1663859327
transform 1 0 40992 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_13_357
timestamp 1663859327
transform 1 0 41328 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_13_389
timestamp 1663859327
transform 1 0 44912 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_13_405
timestamp 1663859327
transform 1 0 46704 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_13_413
timestamp 1663859327
transform 1 0 47600 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_13_417
timestamp 1663859327
transform 1 0 48048 0 -1 14112
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_13_419
timestamp 1663859327
transform 1 0 48272 0 -1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_2
timestamp 1663859327
transform 1 0 1568 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_7
timestamp 1663859327
transform 1 0 2128 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_23
timestamp 1663859327
transform 1 0 3920 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_31
timestamp 1663859327
transform 1 0 4816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_37
timestamp 1663859327
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_101
timestamp 1663859327
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_105
timestamp 1663859327
transform 1 0 13104 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_108
timestamp 1663859327
transform 1 0 13440 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_172
timestamp 1663859327
transform 1 0 20608 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_176
timestamp 1663859327
transform 1 0 21056 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_179
timestamp 1663859327
transform 1 0 21392 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_243
timestamp 1663859327
transform 1 0 28560 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_247
timestamp 1663859327
transform 1 0 29008 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_250
timestamp 1663859327
transform 1 0 29344 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_314
timestamp 1663859327
transform 1 0 36512 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_318
timestamp 1663859327
transform 1 0 36960 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_14_321
timestamp 1663859327
transform 1 0 37296 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_385
timestamp 1663859327
transform 1 0 44464 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_14_389
timestamp 1663859327
transform 1 0 44912 0 1 14112
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_14_392
timestamp 1663859327
transform 1 0 45248 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_14_408
timestamp 1663859327
transform 1 0 47040 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_14_416
timestamp 1663859327
transform 1 0 47936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_2
timestamp 1663859327
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_66
timestamp 1663859327
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_70
timestamp 1663859327
transform 1 0 9184 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_73
timestamp 1663859327
transform 1 0 9520 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_137
timestamp 1663859327
transform 1 0 16688 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_141
timestamp 1663859327
transform 1 0 17136 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_144
timestamp 1663859327
transform 1 0 17472 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_208
timestamp 1663859327
transform 1 0 24640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_212
timestamp 1663859327
transform 1 0 25088 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_215
timestamp 1663859327
transform 1 0 25424 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_279
timestamp 1663859327
transform 1 0 32592 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_283
timestamp 1663859327
transform 1 0 33040 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_15_286
timestamp 1663859327
transform 1 0 33376 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_350
timestamp 1663859327
transform 1 0 40544 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_354
timestamp 1663859327
transform 1 0 40992 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_15_357
timestamp 1663859327
transform 1 0 41328 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_15_389
timestamp 1663859327
transform 1 0 44912 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_15_405
timestamp 1663859327
transform 1 0 46704 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_15_413
timestamp 1663859327
transform 1 0 47600 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_15_417
timestamp 1663859327
transform 1 0 48048 0 -1 15680
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_15_419
timestamp 1663859327
transform 1 0 48272 0 -1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_2
timestamp 1663859327
transform 1 0 1568 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_7
timestamp 1663859327
transform 1 0 2128 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_23
timestamp 1663859327
transform 1 0 3920 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_31
timestamp 1663859327
transform 1 0 4816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_37
timestamp 1663859327
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_101
timestamp 1663859327
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_105
timestamp 1663859327
transform 1 0 13104 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_108
timestamp 1663859327
transform 1 0 13440 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_172
timestamp 1663859327
transform 1 0 20608 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_176
timestamp 1663859327
transform 1 0 21056 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_179
timestamp 1663859327
transform 1 0 21392 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_243
timestamp 1663859327
transform 1 0 28560 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_247
timestamp 1663859327
transform 1 0 29008 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_250
timestamp 1663859327
transform 1 0 29344 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_314
timestamp 1663859327
transform 1 0 36512 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_318
timestamp 1663859327
transform 1 0 36960 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_16_321
timestamp 1663859327
transform 1 0 37296 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_385
timestamp 1663859327
transform 1 0 44464 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_16_389
timestamp 1663859327
transform 1 0 44912 0 1 15680
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_16_392
timestamp 1663859327
transform 1 0 45248 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_16_408
timestamp 1663859327
transform 1 0 47040 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_16_416
timestamp 1663859327
transform 1 0 47936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_2
timestamp 1663859327
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_66
timestamp 1663859327
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_70
timestamp 1663859327
transform 1 0 9184 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_73
timestamp 1663859327
transform 1 0 9520 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_137
timestamp 1663859327
transform 1 0 16688 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_141
timestamp 1663859327
transform 1 0 17136 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_144
timestamp 1663859327
transform 1 0 17472 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_208
timestamp 1663859327
transform 1 0 24640 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_212
timestamp 1663859327
transform 1 0 25088 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_215
timestamp 1663859327
transform 1 0 25424 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_279
timestamp 1663859327
transform 1 0 32592 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_283
timestamp 1663859327
transform 1 0 33040 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_17_286
timestamp 1663859327
transform 1 0 33376 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_350
timestamp 1663859327
transform 1 0 40544 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_354
timestamp 1663859327
transform 1 0 40992 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_17_357
timestamp 1663859327
transform 1 0 41328 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_17_389
timestamp 1663859327
transform 1 0 44912 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_17_405
timestamp 1663859327
transform 1 0 46704 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_17_413
timestamp 1663859327
transform 1 0 47600 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_17_417
timestamp 1663859327
transform 1 0 48048 0 -1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_17_419
timestamp 1663859327
transform 1 0 48272 0 -1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_2
timestamp 1663859327
transform 1 0 1568 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_7
timestamp 1663859327
transform 1 0 2128 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_18_23
timestamp 1663859327
transform 1 0 3920 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_31
timestamp 1663859327
transform 1 0 4816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_37
timestamp 1663859327
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_101
timestamp 1663859327
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_105
timestamp 1663859327
transform 1 0 13104 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_108
timestamp 1663859327
transform 1 0 13440 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_172
timestamp 1663859327
transform 1 0 20608 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_176
timestamp 1663859327
transform 1 0 21056 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_179
timestamp 1663859327
transform 1 0 21392 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_243
timestamp 1663859327
transform 1 0 28560 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_247
timestamp 1663859327
transform 1 0 29008 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_250
timestamp 1663859327
transform 1 0 29344 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_314
timestamp 1663859327
transform 1 0 36512 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_318
timestamp 1663859327
transform 1 0 36960 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_18_321
timestamp 1663859327
transform 1 0 37296 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_385
timestamp 1663859327
transform 1 0 44464 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_389
timestamp 1663859327
transform 1 0 44912 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_18_392
timestamp 1663859327
transform 1 0 45248 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_18_408
timestamp 1663859327
transform 1 0 47040 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_18_412
timestamp 1663859327
transform 1 0 47488 0 1 17248
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_414
timestamp 1663859327
transform 1 0 47712 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_18_419
timestamp 1663859327
transform 1 0 48272 0 1 17248
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_2
timestamp 1663859327
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_66
timestamp 1663859327
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_70
timestamp 1663859327
transform 1 0 9184 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_73
timestamp 1663859327
transform 1 0 9520 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_137
timestamp 1663859327
transform 1 0 16688 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_141
timestamp 1663859327
transform 1 0 17136 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_144
timestamp 1663859327
transform 1 0 17472 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_208
timestamp 1663859327
transform 1 0 24640 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_212
timestamp 1663859327
transform 1 0 25088 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_215
timestamp 1663859327
transform 1 0 25424 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_279
timestamp 1663859327
transform 1 0 32592 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_283
timestamp 1663859327
transform 1 0 33040 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_19_286
timestamp 1663859327
transform 1 0 33376 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_19_350
timestamp 1663859327
transform 1 0 40544 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_354
timestamp 1663859327
transform 1 0 40992 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_19_357
timestamp 1663859327
transform 1 0 41328 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_19_389
timestamp 1663859327
transform 1 0 44912 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_19_405
timestamp 1663859327
transform 1 0 46704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_19_413
timestamp 1663859327
transform 1 0 47600 0 -1 18816
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_19_419
timestamp 1663859327
transform 1 0 48272 0 -1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_2
timestamp 1663859327
transform 1 0 1568 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_7
timestamp 1663859327
transform 1 0 2128 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_23
timestamp 1663859327
transform 1 0 3920 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_31
timestamp 1663859327
transform 1 0 4816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_37
timestamp 1663859327
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_101
timestamp 1663859327
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_105
timestamp 1663859327
transform 1 0 13104 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_108
timestamp 1663859327
transform 1 0 13440 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_172
timestamp 1663859327
transform 1 0 20608 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_176
timestamp 1663859327
transform 1 0 21056 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_179
timestamp 1663859327
transform 1 0 21392 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_243
timestamp 1663859327
transform 1 0 28560 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_247
timestamp 1663859327
transform 1 0 29008 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_250
timestamp 1663859327
transform 1 0 29344 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_314
timestamp 1663859327
transform 1 0 36512 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_318
timestamp 1663859327
transform 1 0 36960 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_20_321
timestamp 1663859327
transform 1 0 37296 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_385
timestamp 1663859327
transform 1 0 44464 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_20_389
timestamp 1663859327
transform 1 0 44912 0 1 18816
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_20_392
timestamp 1663859327
transform 1 0 45248 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_20_408
timestamp 1663859327
transform 1 0 47040 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_20_416
timestamp 1663859327
transform 1 0 47936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_2
timestamp 1663859327
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_66
timestamp 1663859327
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_70
timestamp 1663859327
transform 1 0 9184 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_73
timestamp 1663859327
transform 1 0 9520 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_137
timestamp 1663859327
transform 1 0 16688 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_141
timestamp 1663859327
transform 1 0 17136 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_144
timestamp 1663859327
transform 1 0 17472 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_208
timestamp 1663859327
transform 1 0 24640 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_212
timestamp 1663859327
transform 1 0 25088 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_215
timestamp 1663859327
transform 1 0 25424 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_279
timestamp 1663859327
transform 1 0 32592 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_283
timestamp 1663859327
transform 1 0 33040 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_21_286
timestamp 1663859327
transform 1 0 33376 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_350
timestamp 1663859327
transform 1 0 40544 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_354
timestamp 1663859327
transform 1 0 40992 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_21_357
timestamp 1663859327
transform 1 0 41328 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_21_389
timestamp 1663859327
transform 1 0 44912 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_21_405
timestamp 1663859327
transform 1 0 46704 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_21_413
timestamp 1663859327
transform 1 0 47600 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_21_417
timestamp 1663859327
transform 1 0 48048 0 -1 20384
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_21_419
timestamp 1663859327
transform 1 0 48272 0 -1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_22_2
timestamp 1663859327
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_34
timestamp 1663859327
transform 1 0 5152 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_37
timestamp 1663859327
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_101
timestamp 1663859327
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_105
timestamp 1663859327
transform 1 0 13104 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_108
timestamp 1663859327
transform 1 0 13440 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_172
timestamp 1663859327
transform 1 0 20608 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_176
timestamp 1663859327
transform 1 0 21056 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_179
timestamp 1663859327
transform 1 0 21392 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_243
timestamp 1663859327
transform 1 0 28560 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_247
timestamp 1663859327
transform 1 0 29008 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_250
timestamp 1663859327
transform 1 0 29344 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_314
timestamp 1663859327
transform 1 0 36512 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_318
timestamp 1663859327
transform 1 0 36960 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_22_321
timestamp 1663859327
transform 1 0 37296 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_385
timestamp 1663859327
transform 1 0 44464 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_22_389
timestamp 1663859327
transform 1 0 44912 0 1 20384
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_22_392
timestamp 1663859327
transform 1 0 45248 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_22_408
timestamp 1663859327
transform 1 0 47040 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_22_416
timestamp 1663859327
transform 1 0 47936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_2
timestamp 1663859327
transform 1 0 1568 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_7
timestamp 1663859327
transform 1 0 2128 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_73
timestamp 1663859327
transform 1 0 9520 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_137
timestamp 1663859327
transform 1 0 16688 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_141
timestamp 1663859327
transform 1 0 17136 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_144
timestamp 1663859327
transform 1 0 17472 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_208
timestamp 1663859327
transform 1 0 24640 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_212
timestamp 1663859327
transform 1 0 25088 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_215
timestamp 1663859327
transform 1 0 25424 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_279
timestamp 1663859327
transform 1 0 32592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_283
timestamp 1663859327
transform 1 0 33040 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_23_286
timestamp 1663859327
transform 1 0 33376 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_350
timestamp 1663859327
transform 1 0 40544 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_354
timestamp 1663859327
transform 1 0 40992 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_23_357
timestamp 1663859327
transform 1 0 41328 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_23_389
timestamp 1663859327
transform 1 0 44912 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_23_405
timestamp 1663859327
transform 1 0 46704 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_23_413
timestamp 1663859327
transform 1 0 47600 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_23_417
timestamp 1663859327
transform 1 0 48048 0 -1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_23_419
timestamp 1663859327
transform 1 0 48272 0 -1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_24_2
timestamp 1663859327
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_34
timestamp 1663859327
transform 1 0 5152 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_37
timestamp 1663859327
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_101
timestamp 1663859327
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_105
timestamp 1663859327
transform 1 0 13104 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_108
timestamp 1663859327
transform 1 0 13440 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_172
timestamp 1663859327
transform 1 0 20608 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_176
timestamp 1663859327
transform 1 0 21056 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_179
timestamp 1663859327
transform 1 0 21392 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_243
timestamp 1663859327
transform 1 0 28560 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_247
timestamp 1663859327
transform 1 0 29008 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_250
timestamp 1663859327
transform 1 0 29344 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_314
timestamp 1663859327
transform 1 0 36512 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_318
timestamp 1663859327
transform 1 0 36960 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_24_321
timestamp 1663859327
transform 1 0 37296 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_385
timestamp 1663859327
transform 1 0 44464 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_389
timestamp 1663859327
transform 1 0 44912 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_24_392
timestamp 1663859327
transform 1 0 45248 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_24_408
timestamp 1663859327
transform 1 0 47040 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_24_412
timestamp 1663859327
transform 1 0 47488 0 1 21952
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_414
timestamp 1663859327
transform 1 0 47712 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_24_419
timestamp 1663859327
transform 1 0 48272 0 1 21952
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_2
timestamp 1663859327
transform 1 0 1568 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_17
timestamp 1663859327
transform 1 0 3248 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_21
timestamp 1663859327
transform 1 0 3696 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_53
timestamp 1663859327
transform 1 0 7280 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_69
timestamp 1663859327
transform 1 0 9072 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_73
timestamp 1663859327
transform 1 0 9520 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_137
timestamp 1663859327
transform 1 0 16688 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_141
timestamp 1663859327
transform 1 0 17136 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_144
timestamp 1663859327
transform 1 0 17472 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_208
timestamp 1663859327
transform 1 0 24640 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_212
timestamp 1663859327
transform 1 0 25088 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_215
timestamp 1663859327
transform 1 0 25424 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_279
timestamp 1663859327
transform 1 0 32592 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_283
timestamp 1663859327
transform 1 0 33040 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_25_286
timestamp 1663859327
transform 1 0 33376 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_350
timestamp 1663859327
transform 1 0 40544 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_354
timestamp 1663859327
transform 1 0 40992 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_25_357
timestamp 1663859327
transform 1 0 41328 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_25_389
timestamp 1663859327
transform 1 0 44912 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_25_405
timestamp 1663859327
transform 1 0 46704 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_25_413
timestamp 1663859327
transform 1 0 47600 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_25_417
timestamp 1663859327
transform 1 0 48048 0 -1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_25_419
timestamp 1663859327
transform 1 0 48272 0 -1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_26_2
timestamp 1663859327
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_34
timestamp 1663859327
transform 1 0 5152 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_37
timestamp 1663859327
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_101
timestamp 1663859327
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_105
timestamp 1663859327
transform 1 0 13104 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_108
timestamp 1663859327
transform 1 0 13440 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_172
timestamp 1663859327
transform 1 0 20608 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_176
timestamp 1663859327
transform 1 0 21056 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_179
timestamp 1663859327
transform 1 0 21392 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_243
timestamp 1663859327
transform 1 0 28560 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_247
timestamp 1663859327
transform 1 0 29008 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_250
timestamp 1663859327
transform 1 0 29344 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_314
timestamp 1663859327
transform 1 0 36512 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_318
timestamp 1663859327
transform 1 0 36960 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_26_321
timestamp 1663859327
transform 1 0 37296 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_385
timestamp 1663859327
transform 1 0 44464 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_389
timestamp 1663859327
transform 1 0 44912 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_26_392
timestamp 1663859327
transform 1 0 45248 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_26_408
timestamp 1663859327
transform 1 0 47040 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_26_412
timestamp 1663859327
transform 1 0 47488 0 1 23520
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_414
timestamp 1663859327
transform 1 0 47712 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_26_419
timestamp 1663859327
transform 1 0 48272 0 1 23520
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_2
timestamp 1663859327
transform 1 0 1568 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_7
timestamp 1663859327
transform 1 0 2128 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_73
timestamp 1663859327
transform 1 0 9520 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_137
timestamp 1663859327
transform 1 0 16688 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_141
timestamp 1663859327
transform 1 0 17136 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_144
timestamp 1663859327
transform 1 0 17472 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_208
timestamp 1663859327
transform 1 0 24640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_212
timestamp 1663859327
transform 1 0 25088 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_215
timestamp 1663859327
transform 1 0 25424 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_279
timestamp 1663859327
transform 1 0 32592 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_283
timestamp 1663859327
transform 1 0 33040 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_27_286
timestamp 1663859327
transform 1 0 33376 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_350
timestamp 1663859327
transform 1 0 40544 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_354
timestamp 1663859327
transform 1 0 40992 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_27_357
timestamp 1663859327
transform 1 0 41328 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_27_389
timestamp 1663859327
transform 1 0 44912 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_27_405
timestamp 1663859327
transform 1 0 46704 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_27_413
timestamp 1663859327
transform 1 0 47600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_27_417
timestamp 1663859327
transform 1 0 48048 0 -1 25088
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_27_419
timestamp 1663859327
transform 1 0 48272 0 -1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_28_2
timestamp 1663859327
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_34
timestamp 1663859327
transform 1 0 5152 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_37
timestamp 1663859327
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_101
timestamp 1663859327
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_105
timestamp 1663859327
transform 1 0 13104 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_108
timestamp 1663859327
transform 1 0 13440 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_172
timestamp 1663859327
transform 1 0 20608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_176
timestamp 1663859327
transform 1 0 21056 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_179
timestamp 1663859327
transform 1 0 21392 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_243
timestamp 1663859327
transform 1 0 28560 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_247
timestamp 1663859327
transform 1 0 29008 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_250
timestamp 1663859327
transform 1 0 29344 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_314
timestamp 1663859327
transform 1 0 36512 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_318
timestamp 1663859327
transform 1 0 36960 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_28_321
timestamp 1663859327
transform 1 0 37296 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_385
timestamp 1663859327
transform 1 0 44464 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_28_389
timestamp 1663859327
transform 1 0 44912 0 1 25088
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_28_392
timestamp 1663859327
transform 1 0 45248 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_28_408
timestamp 1663859327
transform 1 0 47040 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_28_416
timestamp 1663859327
transform 1 0 47936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_2
timestamp 1663859327
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_66
timestamp 1663859327
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_70
timestamp 1663859327
transform 1 0 9184 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_73
timestamp 1663859327
transform 1 0 9520 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_137
timestamp 1663859327
transform 1 0 16688 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_141
timestamp 1663859327
transform 1 0 17136 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_144
timestamp 1663859327
transform 1 0 17472 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_208
timestamp 1663859327
transform 1 0 24640 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_212
timestamp 1663859327
transform 1 0 25088 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_215
timestamp 1663859327
transform 1 0 25424 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_279
timestamp 1663859327
transform 1 0 32592 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_283
timestamp 1663859327
transform 1 0 33040 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_29_286
timestamp 1663859327
transform 1 0 33376 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_350
timestamp 1663859327
transform 1 0 40544 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_354
timestamp 1663859327
transform 1 0 40992 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_29_357
timestamp 1663859327
transform 1 0 41328 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_29_389
timestamp 1663859327
transform 1 0 44912 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_29_405
timestamp 1663859327
transform 1 0 46704 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_29_413
timestamp 1663859327
transform 1 0 47600 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_29_417
timestamp 1663859327
transform 1 0 48048 0 -1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_29_419
timestamp 1663859327
transform 1 0 48272 0 -1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_2
timestamp 1663859327
transform 1 0 1568 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_7
timestamp 1663859327
transform 1 0 2128 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_30_23
timestamp 1663859327
transform 1 0 3920 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_31
timestamp 1663859327
transform 1 0 4816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_37
timestamp 1663859327
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_101
timestamp 1663859327
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_105
timestamp 1663859327
transform 1 0 13104 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_108
timestamp 1663859327
transform 1 0 13440 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_172
timestamp 1663859327
transform 1 0 20608 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_176
timestamp 1663859327
transform 1 0 21056 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_179
timestamp 1663859327
transform 1 0 21392 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_243
timestamp 1663859327
transform 1 0 28560 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_247
timestamp 1663859327
transform 1 0 29008 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_250
timestamp 1663859327
transform 1 0 29344 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_314
timestamp 1663859327
transform 1 0 36512 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_318
timestamp 1663859327
transform 1 0 36960 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_30_321
timestamp 1663859327
transform 1 0 37296 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_385
timestamp 1663859327
transform 1 0 44464 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_389
timestamp 1663859327
transform 1 0 44912 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_30_392
timestamp 1663859327
transform 1 0 45248 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_30_408
timestamp 1663859327
transform 1 0 47040 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_30_412
timestamp 1663859327
transform 1 0 47488 0 1 26656
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_414
timestamp 1663859327
transform 1 0 47712 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_30_419
timestamp 1663859327
transform 1 0 48272 0 1 26656
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_2
timestamp 1663859327
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_66
timestamp 1663859327
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_70
timestamp 1663859327
transform 1 0 9184 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_73
timestamp 1663859327
transform 1 0 9520 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_137
timestamp 1663859327
transform 1 0 16688 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_141
timestamp 1663859327
transform 1 0 17136 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_144
timestamp 1663859327
transform 1 0 17472 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_208
timestamp 1663859327
transform 1 0 24640 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_212
timestamp 1663859327
transform 1 0 25088 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_215
timestamp 1663859327
transform 1 0 25424 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_279
timestamp 1663859327
transform 1 0 32592 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_283
timestamp 1663859327
transform 1 0 33040 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_31_286
timestamp 1663859327
transform 1 0 33376 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_350
timestamp 1663859327
transform 1 0 40544 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_354
timestamp 1663859327
transform 1 0 40992 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_31_357
timestamp 1663859327
transform 1 0 41328 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_31_389
timestamp 1663859327
transform 1 0 44912 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_31_405
timestamp 1663859327
transform 1 0 46704 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_31_413
timestamp 1663859327
transform 1 0 47600 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_31_417
timestamp 1663859327
transform 1 0 48048 0 -1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_31_419
timestamp 1663859327
transform 1 0 48272 0 -1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_2
timestamp 1663859327
transform 1 0 1568 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_7
timestamp 1663859327
transform 1 0 2128 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_23
timestamp 1663859327
transform 1 0 3920 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_31
timestamp 1663859327
transform 1 0 4816 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_37
timestamp 1663859327
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_101
timestamp 1663859327
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_105
timestamp 1663859327
transform 1 0 13104 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_108
timestamp 1663859327
transform 1 0 13440 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_172
timestamp 1663859327
transform 1 0 20608 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_176
timestamp 1663859327
transform 1 0 21056 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_179
timestamp 1663859327
transform 1 0 21392 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_185
timestamp 1663859327
transform 1 0 22064 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_187
timestamp 1663859327
transform 1 0 22288 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_190
timestamp 1663859327
transform 1 0 22624 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_32_194
timestamp 1663859327
transform 1 0 23072 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_226
timestamp 1663859327
transform 1 0 26656 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_242
timestamp 1663859327
transform 1 0 28448 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_32_246
timestamp 1663859327
transform 1 0 28896 0 1 28224
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_250
timestamp 1663859327
transform 1 0 29344 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_314
timestamp 1663859327
transform 1 0 36512 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_318
timestamp 1663859327
transform 1 0 36960 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_32_321
timestamp 1663859327
transform 1 0 37296 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_385
timestamp 1663859327
transform 1 0 44464 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_32_389
timestamp 1663859327
transform 1 0 44912 0 1 28224
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_32_392
timestamp 1663859327
transform 1 0 45248 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_32_408
timestamp 1663859327
transform 1 0 47040 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_32_416
timestamp 1663859327
transform 1 0 47936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_2
timestamp 1663859327
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_66
timestamp 1663859327
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_70
timestamp 1663859327
transform 1 0 9184 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_73
timestamp 1663859327
transform 1 0 9520 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_137
timestamp 1663859327
transform 1 0 16688 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_141
timestamp 1663859327
transform 1 0 17136 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_144
timestamp 1663859327
transform 1 0 17472 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_152
timestamp 1663859327
transform 1 0 18368 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_156
timestamp 1663859327
transform 1 0 18816 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_160
timestamp 1663859327
transform 1 0 19264 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_166
timestamp 1663859327
transform 1 0 19936 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_170
timestamp 1663859327
transform 1 0 20384 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_174
timestamp 1663859327
transform 1 0 20832 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_178
timestamp 1663859327
transform 1 0 21280 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_182
timestamp 1663859327
transform 1 0 21728 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_186
timestamp 1663859327
transform 1 0 22176 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_190
timestamp 1663859327
transform 1 0 22624 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_194
timestamp 1663859327
transform 1 0 23072 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_198
timestamp 1663859327
transform 1 0 23520 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_202
timestamp 1663859327
transform 1 0 23968 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_210
timestamp 1663859327
transform 1 0 24864 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_212
timestamp 1663859327
transform 1 0 25088 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_215
timestamp 1663859327
transform 1 0 25424 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_279
timestamp 1663859327
transform 1 0 32592 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_283
timestamp 1663859327
transform 1 0 33040 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_33_286
timestamp 1663859327
transform 1 0 33376 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_33_350
timestamp 1663859327
transform 1 0 40544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_354
timestamp 1663859327
transform 1 0 40992 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_33_357
timestamp 1663859327
transform 1 0 41328 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_33_389
timestamp 1663859327
transform 1 0 44912 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_33_405
timestamp 1663859327
transform 1 0 46704 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_33_413
timestamp 1663859327
transform 1 0 47600 0 -1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_33_419
timestamp 1663859327
transform 1 0 48272 0 -1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_2
timestamp 1663859327
transform 1 0 1568 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_7
timestamp 1663859327
transform 1 0 2128 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_23
timestamp 1663859327
transform 1 0 3920 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_31
timestamp 1663859327
transform 1 0 4816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_37
timestamp 1663859327
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_101
timestamp 1663859327
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_105
timestamp 1663859327
transform 1 0 13104 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_108
timestamp 1663859327
transform 1 0 13440 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_124
timestamp 1663859327
transform 1 0 15232 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_128
timestamp 1663859327
transform 1 0 15680 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_130
timestamp 1663859327
transform 1 0 15904 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_133
timestamp 1663859327
transform 1 0 16240 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_143
timestamp 1663859327
transform 1 0 17360 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_145
timestamp 1663859327
transform 1 0 17584 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_148
timestamp 1663859327
transform 1 0 17920 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_152
timestamp 1663859327
transform 1 0 18368 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_156
timestamp 1663859327
transform 1 0 18816 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_160
timestamp 1663859327
transform 1 0 19264 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_164
timestamp 1663859327
transform 1 0 19712 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_168
timestamp 1663859327
transform 1 0 20160 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_176
timestamp 1663859327
transform 1 0 21056 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_179
timestamp 1663859327
transform 1 0 21392 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_186
timestamp 1663859327
transform 1 0 22176 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_190
timestamp 1663859327
transform 1 0 22624 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_194
timestamp 1663859327
transform 1 0 23072 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_198
timestamp 1663859327
transform 1 0 23520 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_202
timestamp 1663859327
transform 1 0 23968 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_206
timestamp 1663859327
transform 1 0 24416 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_210
timestamp 1663859327
transform 1 0 24864 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_34_214
timestamp 1663859327
transform 1 0 25312 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_34_246
timestamp 1663859327
transform 1 0 28896 0 1 29792
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_250
timestamp 1663859327
transform 1 0 29344 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_314
timestamp 1663859327
transform 1 0 36512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_318
timestamp 1663859327
transform 1 0 36960 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_34_321
timestamp 1663859327
transform 1 0 37296 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_385
timestamp 1663859327
transform 1 0 44464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_34_389
timestamp 1663859327
transform 1 0 44912 0 1 29792
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_34_392
timestamp 1663859327
transform 1 0 45248 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_34_408
timestamp 1663859327
transform 1 0 47040 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_34_416
timestamp 1663859327
transform 1 0 47936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_2
timestamp 1663859327
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_66
timestamp 1663859327
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_70
timestamp 1663859327
transform 1 0 9184 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_73
timestamp 1663859327
transform 1 0 9520 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_105
timestamp 1663859327
transform 1 0 13104 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_113
timestamp 1663859327
transform 1 0 14000 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_117
timestamp 1663859327
transform 1 0 14448 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_121
timestamp 1663859327
transform 1 0 14896 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_125
timestamp 1663859327
transform 1 0 15344 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_129
timestamp 1663859327
transform 1 0 15792 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_133
timestamp 1663859327
transform 1 0 16240 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_137
timestamp 1663859327
transform 1 0 16688 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_141
timestamp 1663859327
transform 1 0 17136 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_144
timestamp 1663859327
transform 1 0 17472 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_147
timestamp 1663859327
transform 1 0 17808 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_151
timestamp 1663859327
transform 1 0 18256 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_155
timestamp 1663859327
transform 1 0 18704 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_159
timestamp 1663859327
transform 1 0 19152 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_167
timestamp 1663859327
transform 1 0 20048 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_177
timestamp 1663859327
transform 1 0 21168 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_187
timestamp 1663859327
transform 1 0 22288 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_195
timestamp 1663859327
transform 1 0 23184 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_199
timestamp 1663859327
transform 1 0 23632 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_203
timestamp 1663859327
transform 1 0 24080 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_207
timestamp 1663859327
transform 1 0 24528 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_211
timestamp 1663859327
transform 1 0 24976 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_215
timestamp 1663859327
transform 1 0 25424 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_218
timestamp 1663859327
transform 1 0 25760 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_222
timestamp 1663859327
transform 1 0 26208 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_254
timestamp 1663859327
transform 1 0 29792 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_270
timestamp 1663859327
transform 1 0 31584 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_278
timestamp 1663859327
transform 1 0 32480 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_282
timestamp 1663859327
transform 1 0 32928 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_35_286
timestamp 1663859327
transform 1 0 33376 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_350
timestamp 1663859327
transform 1 0 40544 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_354
timestamp 1663859327
transform 1 0 40992 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_35_357
timestamp 1663859327
transform 1 0 41328 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_35_389
timestamp 1663859327
transform 1 0 44912 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_35_405
timestamp 1663859327
transform 1 0 46704 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_35_413
timestamp 1663859327
transform 1 0 47600 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_35_417
timestamp 1663859327
transform 1 0 48048 0 -1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_35_419
timestamp 1663859327
transform 1 0 48272 0 -1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_36_2
timestamp 1663859327
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_34
timestamp 1663859327
transform 1 0 5152 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_37
timestamp 1663859327
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_101
timestamp 1663859327
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_105
timestamp 1663859327
transform 1 0 13104 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_108
timestamp 1663859327
transform 1 0 13440 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_112
timestamp 1663859327
transform 1 0 13888 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_116
timestamp 1663859327
transform 1 0 14336 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_120
timestamp 1663859327
transform 1 0 14784 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_124
timestamp 1663859327
transform 1 0 15232 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_128
timestamp 1663859327
transform 1 0 15680 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_132
timestamp 1663859327
transform 1 0 16128 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_136
timestamp 1663859327
transform 1 0 16576 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_140
timestamp 1663859327
transform 1 0 17024 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_144
timestamp 1663859327
transform 1 0 17472 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_148
timestamp 1663859327
transform 1 0 17920 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_156
timestamp 1663859327
transform 1 0 18816 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_164
timestamp 1663859327
transform 1 0 19712 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_176
timestamp 1663859327
transform 1 0 21056 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_179
timestamp 1663859327
transform 1 0 21392 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_188
timestamp 1663859327
transform 1 0 22400 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_197
timestamp 1663859327
transform 1 0 23408 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_205
timestamp 1663859327
transform 1 0 24304 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_209
timestamp 1663859327
transform 1 0 24752 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_211
timestamp 1663859327
transform 1 0 24976 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_214
timestamp 1663859327
transform 1 0 25312 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_218
timestamp 1663859327
transform 1 0 25760 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_222
timestamp 1663859327
transform 1 0 26208 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_226
timestamp 1663859327
transform 1 0 26656 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_230
timestamp 1663859327
transform 1 0 27104 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_246
timestamp 1663859327
transform 1 0 28896 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_250
timestamp 1663859327
transform 1 0 29344 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_314
timestamp 1663859327
transform 1 0 36512 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_318
timestamp 1663859327
transform 1 0 36960 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_36_321
timestamp 1663859327
transform 1 0 37296 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_385
timestamp 1663859327
transform 1 0 44464 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_389
timestamp 1663859327
transform 1 0 44912 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_36_392
timestamp 1663859327
transform 1 0 45248 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_36_408
timestamp 1663859327
transform 1 0 47040 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_36_412
timestamp 1663859327
transform 1 0 47488 0 1 31360
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_414
timestamp 1663859327
transform 1 0 47712 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_36_419
timestamp 1663859327
transform 1 0 48272 0 1 31360
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_2
timestamp 1663859327
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_66
timestamp 1663859327
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_70
timestamp 1663859327
transform 1 0 9184 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_73
timestamp 1663859327
transform 1 0 9520 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_89
timestamp 1663859327
transform 1 0 11312 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_93
timestamp 1663859327
transform 1 0 11760 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_95
timestamp 1663859327
transform 1 0 11984 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_98
timestamp 1663859327
transform 1 0 12320 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_102
timestamp 1663859327
transform 1 0 12768 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_106
timestamp 1663859327
transform 1 0 13216 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_110
timestamp 1663859327
transform 1 0 13664 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_114
timestamp 1663859327
transform 1 0 14112 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_118
timestamp 1663859327
transform 1 0 14560 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_122
timestamp 1663859327
transform 1 0 15008 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_126
timestamp 1663859327
transform 1 0 15456 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_130
timestamp 1663859327
transform 1 0 15904 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_134
timestamp 1663859327
transform 1 0 16352 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_141
timestamp 1663859327
transform 1 0 17136 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_144
timestamp 1663859327
transform 1 0 17472 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_148
timestamp 1663859327
transform 1 0 17920 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_158
timestamp 1663859327
transform 1 0 19040 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_170
timestamp 1663859327
transform 1 0 20384 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_183
timestamp 1663859327
transform 1 0 21840 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_195
timestamp 1663859327
transform 1 0 23184 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_204
timestamp 1663859327
transform 1 0 24192 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_212
timestamp 1663859327
transform 1 0 25088 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_215
timestamp 1663859327
transform 1 0 25424 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_218
timestamp 1663859327
transform 1 0 25760 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_222
timestamp 1663859327
transform 1 0 26208 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_226
timestamp 1663859327
transform 1 0 26656 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_230
timestamp 1663859327
transform 1 0 27104 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_234
timestamp 1663859327
transform 1 0 27552 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_238
timestamp 1663859327
transform 1 0 28000 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_242
timestamp 1663859327
transform 1 0 28448 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_274
timestamp 1663859327
transform 1 0 32032 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_282
timestamp 1663859327
transform 1 0 32928 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_37_286
timestamp 1663859327
transform 1 0 33376 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_37_350
timestamp 1663859327
transform 1 0 40544 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_354
timestamp 1663859327
transform 1 0 40992 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_37_357
timestamp 1663859327
transform 1 0 41328 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_37_389
timestamp 1663859327
transform 1 0 44912 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_37_405
timestamp 1663859327
transform 1 0 46704 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_37_413
timestamp 1663859327
transform 1 0 47600 0 -1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_37_419
timestamp 1663859327
transform 1 0 48272 0 -1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_2
timestamp 1663859327
transform 1 0 1568 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_7
timestamp 1663859327
transform 1 0 2128 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_15
timestamp 1663859327
transform 1 0 3024 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_19
timestamp 1663859327
transform 1 0 3472 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_21
timestamp 1663859327
transform 1 0 3696 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_24
timestamp 1663859327
transform 1 0 4032 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_32
timestamp 1663859327
transform 1 0 4928 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_34
timestamp 1663859327
transform 1 0 5152 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_38_37
timestamp 1663859327
transform 1 0 5488 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_69
timestamp 1663859327
transform 1 0 9072 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_87
timestamp 1663859327
transform 1 0 11088 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_93
timestamp 1663859327
transform 1 0 11760 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_97
timestamp 1663859327
transform 1 0 12208 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_101
timestamp 1663859327
transform 1 0 12656 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_105
timestamp 1663859327
transform 1 0 13104 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_108
timestamp 1663859327
transform 1 0 13440 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_111
timestamp 1663859327
transform 1 0 13776 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_115
timestamp 1663859327
transform 1 0 14224 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_119
timestamp 1663859327
transform 1 0 14672 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_123
timestamp 1663859327
transform 1 0 15120 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_127
timestamp 1663859327
transform 1 0 15568 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_131
timestamp 1663859327
transform 1 0 16016 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_139
timestamp 1663859327
transform 1 0 16912 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_147
timestamp 1663859327
transform 1 0 17808 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_157
timestamp 1663859327
transform 1 0 18928 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_172
timestamp 1663859327
transform 1 0 20608 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_176
timestamp 1663859327
transform 1 0 21056 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_179
timestamp 1663859327
transform 1 0 21392 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_192
timestamp 1663859327
transform 1 0 22848 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_204
timestamp 1663859327
transform 1 0 24192 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_212
timestamp 1663859327
transform 1 0 25088 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_220
timestamp 1663859327
transform 1 0 25984 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_226
timestamp 1663859327
transform 1 0 26656 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_230
timestamp 1663859327
transform 1 0 27104 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_234
timestamp 1663859327
transform 1 0 27552 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_238
timestamp 1663859327
transform 1 0 28000 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_242
timestamp 1663859327
transform 1 0 28448 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_246
timestamp 1663859327
transform 1 0 28896 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_250
timestamp 1663859327
transform 1 0 29344 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_253
timestamp 1663859327
transform 1 0 29680 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_38_317
timestamp 1663859327
transform 1 0 36848 0 1 32928
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_38_321
timestamp 1663859327
transform 1 0 37296 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_385
timestamp 1663859327
transform 1 0 44464 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_38_389
timestamp 1663859327
transform 1 0 44912 0 1 32928
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_38_392
timestamp 1663859327
transform 1 0 45248 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_38_408
timestamp 1663859327
transform 1 0 47040 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_38_416
timestamp 1663859327
transform 1 0 47936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_2
timestamp 1663859327
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_66
timestamp 1663859327
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_70
timestamp 1663859327
transform 1 0 9184 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_73
timestamp 1663859327
transform 1 0 9520 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_76
timestamp 1663859327
transform 1 0 9856 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_80
timestamp 1663859327
transform 1 0 10304 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_84
timestamp 1663859327
transform 1 0 10752 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_88
timestamp 1663859327
transform 1 0 11200 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_92
timestamp 1663859327
transform 1 0 11648 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_96
timestamp 1663859327
transform 1 0 12096 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_100
timestamp 1663859327
transform 1 0 12544 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_104
timestamp 1663859327
transform 1 0 12992 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_108
timestamp 1663859327
transform 1 0 13440 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_112
timestamp 1663859327
transform 1 0 13888 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_116
timestamp 1663859327
transform 1 0 14336 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_124
timestamp 1663859327
transform 1 0 15232 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_132
timestamp 1663859327
transform 1 0 16128 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_141
timestamp 1663859327
transform 1 0 17136 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_144
timestamp 1663859327
transform 1 0 17472 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_155
timestamp 1663859327
transform 1 0 18704 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_186
timestamp 1663859327
transform 1 0 22176 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_201
timestamp 1663859327
transform 1 0 23856 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_212
timestamp 1663859327
transform 1 0 25088 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_215
timestamp 1663859327
transform 1 0 25424 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_222
timestamp 1663859327
transform 1 0 26208 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_230
timestamp 1663859327
transform 1 0 27104 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_236
timestamp 1663859327
transform 1 0 27776 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_240
timestamp 1663859327
transform 1 0 28224 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_244
timestamp 1663859327
transform 1 0 28672 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_248
timestamp 1663859327
transform 1 0 29120 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_252
timestamp 1663859327
transform 1 0 29568 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_256
timestamp 1663859327
transform 1 0 30016 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_260
timestamp 1663859327
transform 1 0 30464 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_264
timestamp 1663859327
transform 1 0 30912 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_268
timestamp 1663859327
transform 1 0 31360 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_39_286
timestamp 1663859327
transform 1 0 33376 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_350
timestamp 1663859327
transform 1 0 40544 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_354
timestamp 1663859327
transform 1 0 40992 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_39_357
timestamp 1663859327
transform 1 0 41328 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_39_389
timestamp 1663859327
transform 1 0 44912 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_39_405
timestamp 1663859327
transform 1 0 46704 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_39_413
timestamp 1663859327
transform 1 0 47600 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_39_417
timestamp 1663859327
transform 1 0 48048 0 -1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_39_419
timestamp 1663859327
transform 1 0 48272 0 -1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_2
timestamp 1663859327
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_34
timestamp 1663859327
transform 1 0 5152 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_37
timestamp 1663859327
transform 1 0 5488 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_40_53
timestamp 1663859327
transform 1 0 7280 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_61
timestamp 1663859327
transform 1 0 8176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_65
timestamp 1663859327
transform 1 0 8624 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_69
timestamp 1663859327
transform 1 0 9072 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_73
timestamp 1663859327
transform 1 0 9520 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_77
timestamp 1663859327
transform 1 0 9968 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_81
timestamp 1663859327
transform 1 0 10416 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_85
timestamp 1663859327
transform 1 0 10864 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_89
timestamp 1663859327
transform 1 0 11312 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_93
timestamp 1663859327
transform 1 0 11760 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_97
timestamp 1663859327
transform 1 0 12208 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_101
timestamp 1663859327
transform 1 0 12656 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_105
timestamp 1663859327
transform 1 0 13104 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_108
timestamp 1663859327
transform 1 0 13440 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_116
timestamp 1663859327
transform 1 0 14336 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_124
timestamp 1663859327
transform 1 0 15232 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_133
timestamp 1663859327
transform 1 0 16240 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_145
timestamp 1663859327
transform 1 0 17584 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_176
timestamp 1663859327
transform 1 0 21056 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_179
timestamp 1663859327
transform 1 0 21392 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_209
timestamp 1663859327
transform 1 0 24752 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_221
timestamp 1663859327
transform 1 0 26096 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_231
timestamp 1663859327
transform 1 0 27216 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_239
timestamp 1663859327
transform 1 0 28112 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_245
timestamp 1663859327
transform 1 0 28784 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_247
timestamp 1663859327
transform 1 0 29008 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_250
timestamp 1663859327
transform 1 0 29344 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_253
timestamp 1663859327
transform 1 0 29680 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_257
timestamp 1663859327
transform 1 0 30128 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_261
timestamp 1663859327
transform 1 0 30576 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_265
timestamp 1663859327
transform 1 0 31024 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_269
timestamp 1663859327
transform 1 0 31472 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_273
timestamp 1663859327
transform 1 0 31920 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_277
timestamp 1663859327
transform 1 0 32368 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_40_281
timestamp 1663859327
transform 1 0 32816 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_313
timestamp 1663859327
transform 1 0 36400 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_317
timestamp 1663859327
transform 1 0 36848 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_40_321
timestamp 1663859327
transform 1 0 37296 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_385
timestamp 1663859327
transform 1 0 44464 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_389
timestamp 1663859327
transform 1 0 44912 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_40_392
timestamp 1663859327
transform 1 0 45248 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_40_408
timestamp 1663859327
transform 1 0 47040 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_40_412
timestamp 1663859327
transform 1 0 47488 0 1 34496
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_414
timestamp 1663859327
transform 1 0 47712 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_40_419
timestamp 1663859327
transform 1 0 48272 0 1 34496
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_2
timestamp 1663859327
transform 1 0 1568 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_7
timestamp 1663859327
transform 1 0 2128 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_39
timestamp 1663859327
transform 1 0 5712 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_47
timestamp 1663859327
transform 1 0 6608 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_51
timestamp 1663859327
transform 1 0 7056 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_54
timestamp 1663859327
transform 1 0 7392 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_58
timestamp 1663859327
transform 1 0 7840 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_62
timestamp 1663859327
transform 1 0 8288 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_66
timestamp 1663859327
transform 1 0 8736 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_70
timestamp 1663859327
transform 1 0 9184 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_73
timestamp 1663859327
transform 1 0 9520 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_77
timestamp 1663859327
transform 1 0 9968 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_81
timestamp 1663859327
transform 1 0 10416 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_85
timestamp 1663859327
transform 1 0 10864 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_89
timestamp 1663859327
transform 1 0 11312 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_93
timestamp 1663859327
transform 1 0 11760 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_97
timestamp 1663859327
transform 1 0 12208 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_103
timestamp 1663859327
transform 1 0 12880 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_111
timestamp 1663859327
transform 1 0 13776 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_119
timestamp 1663859327
transform 1 0 14672 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_129
timestamp 1663859327
transform 1 0 15792 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_141
timestamp 1663859327
transform 1 0 17136 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_144
timestamp 1663859327
transform 1 0 17472 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_157
timestamp 1663859327
transform 1 0 18928 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_188
timestamp 1663859327
transform 1 0 22400 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_206
timestamp 1663859327
transform 1 0 24416 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_212
timestamp 1663859327
transform 1 0 25088 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_215
timestamp 1663859327
transform 1 0 25424 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_227
timestamp 1663859327
transform 1 0 26768 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_237
timestamp 1663859327
transform 1 0 27888 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_245
timestamp 1663859327
transform 1 0 28784 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_251
timestamp 1663859327
transform 1 0 29456 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_255
timestamp 1663859327
transform 1 0 29904 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_259
timestamp 1663859327
transform 1 0 30352 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_263
timestamp 1663859327
transform 1 0 30800 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_267
timestamp 1663859327
transform 1 0 31248 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_271
timestamp 1663859327
transform 1 0 31696 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_275
timestamp 1663859327
transform 1 0 32144 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_279
timestamp 1663859327
transform 1 0 32592 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_283
timestamp 1663859327
transform 1 0 33040 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_286
timestamp 1663859327
transform 1 0 33376 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_41_289
timestamp 1663859327
transform 1 0 33712 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_353
timestamp 1663859327
transform 1 0 40880 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_41_357
timestamp 1663859327
transform 1 0 41328 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_41_389
timestamp 1663859327
transform 1 0 44912 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_41_405
timestamp 1663859327
transform 1 0 46704 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_41_413
timestamp 1663859327
transform 1 0 47600 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_41_417
timestamp 1663859327
transform 1 0 48048 0 -1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_41_419
timestamp 1663859327
transform 1 0 48272 0 -1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_42_2
timestamp 1663859327
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_34
timestamp 1663859327
transform 1 0 5152 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_37
timestamp 1663859327
transform 1 0 5488 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_41
timestamp 1663859327
transform 1 0 5936 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_45
timestamp 1663859327
transform 1 0 6384 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_49
timestamp 1663859327
transform 1 0 6832 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_53
timestamp 1663859327
transform 1 0 7280 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_57
timestamp 1663859327
transform 1 0 7728 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_61
timestamp 1663859327
transform 1 0 8176 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_65
timestamp 1663859327
transform 1 0 8624 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_69
timestamp 1663859327
transform 1 0 9072 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_73
timestamp 1663859327
transform 1 0 9520 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_77
timestamp 1663859327
transform 1 0 9968 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_81
timestamp 1663859327
transform 1 0 10416 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_85
timestamp 1663859327
transform 1 0 10864 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_89
timestamp 1663859327
transform 1 0 11312 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_97
timestamp 1663859327
transform 1 0 12208 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_105
timestamp 1663859327
transform 1 0 13104 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_108
timestamp 1663859327
transform 1 0 13440 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_114
timestamp 1663859327
transform 1 0 14112 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_145
timestamp 1663859327
transform 1 0 17584 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_176
timestamp 1663859327
transform 1 0 21056 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_179
timestamp 1663859327
transform 1 0 21392 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_209
timestamp 1663859327
transform 1 0 24752 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_224
timestamp 1663859327
transform 1 0 26432 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_237
timestamp 1663859327
transform 1 0 27888 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_247
timestamp 1663859327
transform 1 0 29008 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_250
timestamp 1663859327
transform 1 0 29344 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_257
timestamp 1663859327
transform 1 0 30128 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_261
timestamp 1663859327
transform 1 0 30576 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_265
timestamp 1663859327
transform 1 0 31024 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_269
timestamp 1663859327
transform 1 0 31472 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_273
timestamp 1663859327
transform 1 0 31920 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_277
timestamp 1663859327
transform 1 0 32368 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_281
timestamp 1663859327
transform 1 0 32816 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_285
timestamp 1663859327
transform 1 0 33264 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_289
timestamp 1663859327
transform 1 0 33712 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_293
timestamp 1663859327
transform 1 0 34160 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_297
timestamp 1663859327
transform 1 0 34608 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_301
timestamp 1663859327
transform 1 0 35056 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_317
timestamp 1663859327
transform 1 0 36848 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_42_321
timestamp 1663859327
transform 1 0 37296 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_385
timestamp 1663859327
transform 1 0 44464 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_389
timestamp 1663859327
transform 1 0 44912 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_42_392
timestamp 1663859327
transform 1 0 45248 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_42_408
timestamp 1663859327
transform 1 0 47040 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_42_412
timestamp 1663859327
transform 1 0 47488 0 1 36064
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_414
timestamp 1663859327
transform 1 0 47712 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_42_419
timestamp 1663859327
transform 1 0 48272 0 1 36064
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_2
timestamp 1663859327
transform 1 0 1568 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_7
timestamp 1663859327
transform 1 0 2128 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_23
timestamp 1663859327
transform 1 0 3920 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_31
timestamp 1663859327
transform 1 0 4816 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_35
timestamp 1663859327
transform 1 0 5264 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_38
timestamp 1663859327
transform 1 0 5600 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_42
timestamp 1663859327
transform 1 0 6048 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_46
timestamp 1663859327
transform 1 0 6496 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_50
timestamp 1663859327
transform 1 0 6944 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_54
timestamp 1663859327
transform 1 0 7392 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_58
timestamp 1663859327
transform 1 0 7840 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_62
timestamp 1663859327
transform 1 0 8288 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_66
timestamp 1663859327
transform 1 0 8736 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_70
timestamp 1663859327
transform 1 0 9184 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_73
timestamp 1663859327
transform 1 0 9520 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_75
timestamp 1663859327
transform 1 0 9744 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_78
timestamp 1663859327
transform 1 0 10080 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_84
timestamp 1663859327
transform 1 0 10752 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_92
timestamp 1663859327
transform 1 0 11648 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_100
timestamp 1663859327
transform 1 0 12544 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_110
timestamp 1663859327
transform 1 0 13664 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_141
timestamp 1663859327
transform 1 0 17136 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_144
timestamp 1663859327
transform 1 0 17472 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_159
timestamp 1663859327
transform 1 0 19152 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_190
timestamp 1663859327
transform 1 0 22624 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_209
timestamp 1663859327
transform 1 0 24752 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_215
timestamp 1663859327
transform 1 0 25424 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_239
timestamp 1663859327
transform 1 0 28112 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_251
timestamp 1663859327
transform 1 0 29456 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_261
timestamp 1663859327
transform 1 0 30576 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_269
timestamp 1663859327
transform 1 0 31472 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_273
timestamp 1663859327
transform 1 0 31920 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_277
timestamp 1663859327
transform 1 0 32368 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_281
timestamp 1663859327
transform 1 0 32816 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_283
timestamp 1663859327
transform 1 0 33040 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_286
timestamp 1663859327
transform 1 0 33376 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_289
timestamp 1663859327
transform 1 0 33712 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_293
timestamp 1663859327
transform 1 0 34160 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_297
timestamp 1663859327
transform 1 0 34608 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_301
timestamp 1663859327
transform 1 0 35056 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_305
timestamp 1663859327
transform 1 0 35504 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_309
timestamp 1663859327
transform 1 0 35952 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_341
timestamp 1663859327
transform 1 0 39536 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_349
timestamp 1663859327
transform 1 0 40432 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_353
timestamp 1663859327
transform 1 0 40880 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_43_357
timestamp 1663859327
transform 1 0 41328 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_43_389
timestamp 1663859327
transform 1 0 44912 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_43_405
timestamp 1663859327
transform 1 0 46704 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_43_413
timestamp 1663859327
transform 1 0 47600 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_43_417
timestamp 1663859327
transform 1 0 48048 0 -1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_43_419
timestamp 1663859327
transform 1 0 48272 0 -1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_2
timestamp 1663859327
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_18
timestamp 1663859327
transform 1 0 3360 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_22
timestamp 1663859327
transform 1 0 3808 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_26
timestamp 1663859327
transform 1 0 4256 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_30
timestamp 1663859327
transform 1 0 4704 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_34
timestamp 1663859327
transform 1 0 5152 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_37
timestamp 1663859327
transform 1 0 5488 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_41
timestamp 1663859327
transform 1 0 5936 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_45
timestamp 1663859327
transform 1 0 6384 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_49
timestamp 1663859327
transform 1 0 6832 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_53
timestamp 1663859327
transform 1 0 7280 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_57
timestamp 1663859327
transform 1 0 7728 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_61
timestamp 1663859327
transform 1 0 8176 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_65
timestamp 1663859327
transform 1 0 8624 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_69
timestamp 1663859327
transform 1 0 9072 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_73
timestamp 1663859327
transform 1 0 9520 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_77
timestamp 1663859327
transform 1 0 9968 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_85
timestamp 1663859327
transform 1 0 10864 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_93
timestamp 1663859327
transform 1 0 11760 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_105
timestamp 1663859327
transform 1 0 13104 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_108
timestamp 1663859327
transform 1 0 13440 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_114
timestamp 1663859327
transform 1 0 14112 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_145
timestamp 1663859327
transform 1 0 17584 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_176
timestamp 1663859327
transform 1 0 21056 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_179
timestamp 1663859327
transform 1 0 21392 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_209
timestamp 1663859327
transform 1 0 24752 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_240
timestamp 1663859327
transform 1 0 28224 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_247
timestamp 1663859327
transform 1 0 29008 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_250
timestamp 1663859327
transform 1 0 29344 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_259
timestamp 1663859327
transform 1 0 30352 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_269
timestamp 1663859327
transform 1 0 31472 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_277
timestamp 1663859327
transform 1 0 32368 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_281
timestamp 1663859327
transform 1 0 32816 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_285
timestamp 1663859327
transform 1 0 33264 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_289
timestamp 1663859327
transform 1 0 33712 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_293
timestamp 1663859327
transform 1 0 34160 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_297
timestamp 1663859327
transform 1 0 34608 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_301
timestamp 1663859327
transform 1 0 35056 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_305
timestamp 1663859327
transform 1 0 35504 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_309
timestamp 1663859327
transform 1 0 35952 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_313
timestamp 1663859327
transform 1 0 36400 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_317
timestamp 1663859327
transform 1 0 36848 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_44_321
timestamp 1663859327
transform 1 0 37296 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_385
timestamp 1663859327
transform 1 0 44464 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_389
timestamp 1663859327
transform 1 0 44912 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_44_392
timestamp 1663859327
transform 1 0 45248 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_44_408
timestamp 1663859327
transform 1 0 47040 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_44_412
timestamp 1663859327
transform 1 0 47488 0 1 37632
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_414
timestamp 1663859327
transform 1 0 47712 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_44_419
timestamp 1663859327
transform 1 0 48272 0 1 37632
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_2
timestamp 1663859327
transform 1 0 1568 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_7
timestamp 1663859327
transform 1 0 2128 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_15
timestamp 1663859327
transform 1 0 3024 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_19
timestamp 1663859327
transform 1 0 3472 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_22
timestamp 1663859327
transform 1 0 3808 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_26
timestamp 1663859327
transform 1 0 4256 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_30
timestamp 1663859327
transform 1 0 4704 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_34
timestamp 1663859327
transform 1 0 5152 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_38
timestamp 1663859327
transform 1 0 5600 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_42
timestamp 1663859327
transform 1 0 6048 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_46
timestamp 1663859327
transform 1 0 6496 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_50
timestamp 1663859327
transform 1 0 6944 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_54
timestamp 1663859327
transform 1 0 7392 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_58
timestamp 1663859327
transform 1 0 7840 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_62
timestamp 1663859327
transform 1 0 8288 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_66
timestamp 1663859327
transform 1 0 8736 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_70
timestamp 1663859327
transform 1 0 9184 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_73
timestamp 1663859327
transform 1 0 9520 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_85
timestamp 1663859327
transform 1 0 10864 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_95
timestamp 1663859327
transform 1 0 11984 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_110
timestamp 1663859327
transform 1 0 13664 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_141
timestamp 1663859327
transform 1 0 17136 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_144
timestamp 1663859327
transform 1 0 17472 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_147
timestamp 1663859327
transform 1 0 17808 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_181
timestamp 1663859327
transform 1 0 21616 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_212
timestamp 1663859327
transform 1 0 25088 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_215
timestamp 1663859327
transform 1 0 25424 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_245
timestamp 1663859327
transform 1 0 28784 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_259
timestamp 1663859327
transform 1 0 30352 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_269
timestamp 1663859327
transform 1 0 31472 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_279
timestamp 1663859327
transform 1 0 32592 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_283
timestamp 1663859327
transform 1 0 33040 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_286
timestamp 1663859327
transform 1 0 33376 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_289
timestamp 1663859327
transform 1 0 33712 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_293
timestamp 1663859327
transform 1 0 34160 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_297
timestamp 1663859327
transform 1 0 34608 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_301
timestamp 1663859327
transform 1 0 35056 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_305
timestamp 1663859327
transform 1 0 35504 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_309
timestamp 1663859327
transform 1 0 35952 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_313
timestamp 1663859327
transform 1 0 36400 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_317
timestamp 1663859327
transform 1 0 36848 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_321
timestamp 1663859327
transform 1 0 37296 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_325
timestamp 1663859327
transform 1 0 37744 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_341
timestamp 1663859327
transform 1 0 39536 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_349
timestamp 1663859327
transform 1 0 40432 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_353
timestamp 1663859327
transform 1 0 40880 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_45_357
timestamp 1663859327
transform 1 0 41328 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_45_389
timestamp 1663859327
transform 1 0 44912 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_45_405
timestamp 1663859327
transform 1 0 46704 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_45_413
timestamp 1663859327
transform 1 0 47600 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_45_417
timestamp 1663859327
transform 1 0 48048 0 -1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_45_419
timestamp 1663859327
transform 1 0 48272 0 -1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_2
timestamp 1663859327
transform 1 0 1568 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_5
timestamp 1663859327
transform 1 0 1904 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_7
timestamp 1663859327
transform 1 0 2128 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_10
timestamp 1663859327
transform 1 0 2464 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_14
timestamp 1663859327
transform 1 0 2912 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_18
timestamp 1663859327
transform 1 0 3360 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_22
timestamp 1663859327
transform 1 0 3808 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_26
timestamp 1663859327
transform 1 0 4256 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_30
timestamp 1663859327
transform 1 0 4704 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_34
timestamp 1663859327
transform 1 0 5152 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_37
timestamp 1663859327
transform 1 0 5488 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_40
timestamp 1663859327
transform 1 0 5824 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_44
timestamp 1663859327
transform 1 0 6272 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_48
timestamp 1663859327
transform 1 0 6720 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_52
timestamp 1663859327
transform 1 0 7168 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_56
timestamp 1663859327
transform 1 0 7616 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_64
timestamp 1663859327
transform 1 0 8512 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_74
timestamp 1663859327
transform 1 0 9632 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_105
timestamp 1663859327
transform 1 0 13104 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_108
timestamp 1663859327
transform 1 0 13440 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_114
timestamp 1663859327
transform 1 0 14112 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_145
timestamp 1663859327
transform 1 0 17584 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_176
timestamp 1663859327
transform 1 0 21056 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_179
timestamp 1663859327
transform 1 0 21392 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_209
timestamp 1663859327
transform 1 0 24752 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_240
timestamp 1663859327
transform 1 0 28224 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_247
timestamp 1663859327
transform 1 0 29008 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_250
timestamp 1663859327
transform 1 0 29344 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_263
timestamp 1663859327
transform 1 0 30800 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_275
timestamp 1663859327
transform 1 0 32144 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_285
timestamp 1663859327
transform 1 0 33264 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_293
timestamp 1663859327
transform 1 0 34160 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_299
timestamp 1663859327
transform 1 0 34832 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_303
timestamp 1663859327
transform 1 0 35280 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_307
timestamp 1663859327
transform 1 0 35728 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_311
timestamp 1663859327
transform 1 0 36176 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_315
timestamp 1663859327
transform 1 0 36624 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_46_321
timestamp 1663859327
transform 1 0 37296 0 1 39200
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_324
timestamp 1663859327
transform 1 0 37632 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_328
timestamp 1663859327
transform 1 0 38080 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_332
timestamp 1663859327
transform 1 0 38528 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_46_336
timestamp 1663859327
transform 1 0 38976 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_368
timestamp 1663859327
transform 1 0 42560 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_384
timestamp 1663859327
transform 1 0 44352 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_46_388
timestamp 1663859327
transform 1 0 44800 0 1 39200
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_46_392
timestamp 1663859327
transform 1 0 45248 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_46_408
timestamp 1663859327
transform 1 0 47040 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_46_416
timestamp 1663859327
transform 1 0 47936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_2
timestamp 1663859327
transform 1 0 1568 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_8
timestamp 1663859327
transform 1 0 2240 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_12
timestamp 1663859327
transform 1 0 2688 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_16
timestamp 1663859327
transform 1 0 3136 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_20
timestamp 1663859327
transform 1 0 3584 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_24
timestamp 1663859327
transform 1 0 4032 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_28
timestamp 1663859327
transform 1 0 4480 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_32
timestamp 1663859327
transform 1 0 4928 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_36
timestamp 1663859327
transform 1 0 5376 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_40
timestamp 1663859327
transform 1 0 5824 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_44
timestamp 1663859327
transform 1 0 6272 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_52
timestamp 1663859327
transform 1 0 7168 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_60
timestamp 1663859327
transform 1 0 8064 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_70
timestamp 1663859327
transform 1 0 9184 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_73
timestamp 1663859327
transform 1 0 9520 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_79
timestamp 1663859327
transform 1 0 10192 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_110
timestamp 1663859327
transform 1 0 13664 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_141
timestamp 1663859327
transform 1 0 17136 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_144
timestamp 1663859327
transform 1 0 17472 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_153
timestamp 1663859327
transform 1 0 18480 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_189
timestamp 1663859327
transform 1 0 22512 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_209
timestamp 1663859327
transform 1 0 24752 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_215
timestamp 1663859327
transform 1 0 25424 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_245
timestamp 1663859327
transform 1 0 28784 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_270
timestamp 1663859327
transform 1 0 31584 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_282
timestamp 1663859327
transform 1 0 32928 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_286
timestamp 1663859327
transform 1 0 33376 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_295
timestamp 1663859327
transform 1 0 34384 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_303
timestamp 1663859327
transform 1 0 35280 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_307
timestamp 1663859327
transform 1 0 35728 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_311
timestamp 1663859327
transform 1 0 36176 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_315
timestamp 1663859327
transform 1 0 36624 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_319
timestamp 1663859327
transform 1 0 37072 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_323
timestamp 1663859327
transform 1 0 37520 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_327
timestamp 1663859327
transform 1 0 37968 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_331
timestamp 1663859327
transform 1 0 38416 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_335
timestamp 1663859327
transform 1 0 38864 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_339
timestamp 1663859327
transform 1 0 39312 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_343
timestamp 1663859327
transform 1 0 39760 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_47_351
timestamp 1663859327
transform 1 0 40656 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_47_357
timestamp 1663859327
transform 1 0 41328 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_47_389
timestamp 1663859327
transform 1 0 44912 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_47_405
timestamp 1663859327
transform 1 0 46704 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_47_413
timestamp 1663859327
transform 1 0 47600 0 -1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_47_419
timestamp 1663859327
transform 1 0 48272 0 -1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_2
timestamp 1663859327
transform 1 0 1568 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_6
timestamp 1663859327
transform 1 0 2016 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_10
timestamp 1663859327
transform 1 0 2464 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_14
timestamp 1663859327
transform 1 0 2912 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_18
timestamp 1663859327
transform 1 0 3360 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_22
timestamp 1663859327
transform 1 0 3808 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_26
timestamp 1663859327
transform 1 0 4256 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_30
timestamp 1663859327
transform 1 0 4704 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_34
timestamp 1663859327
transform 1 0 5152 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_37
timestamp 1663859327
transform 1 0 5488 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_44
timestamp 1663859327
transform 1 0 6272 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_52
timestamp 1663859327
transform 1 0 7168 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_62
timestamp 1663859327
transform 1 0 8288 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_74
timestamp 1663859327
transform 1 0 9632 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_105
timestamp 1663859327
transform 1 0 13104 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_108
timestamp 1663859327
transform 1 0 13440 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_134
timestamp 1663859327
transform 1 0 16352 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_170
timestamp 1663859327
transform 1 0 20384 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_176
timestamp 1663859327
transform 1 0 21056 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_179
timestamp 1663859327
transform 1 0 21392 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_223
timestamp 1663859327
transform 1 0 26320 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_242
timestamp 1663859327
transform 1 0 28448 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_246
timestamp 1663859327
transform 1 0 28896 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_250
timestamp 1663859327
transform 1 0 29344 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_280
timestamp 1663859327
transform 1 0 32704 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_292
timestamp 1663859327
transform 1 0 34048 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_302
timestamp 1663859327
transform 1 0 35168 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_310
timestamp 1663859327
transform 1 0 36064 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_318
timestamp 1663859327
transform 1 0 36960 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_48_321
timestamp 1663859327
transform 1 0 37296 0 1 40768
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_324
timestamp 1663859327
transform 1 0 37632 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_328
timestamp 1663859327
transform 1 0 38080 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_332
timestamp 1663859327
transform 1 0 38528 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_336
timestamp 1663859327
transform 1 0 38976 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_340
timestamp 1663859327
transform 1 0 39424 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_344
timestamp 1663859327
transform 1 0 39872 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_348
timestamp 1663859327
transform 1 0 40320 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_48_352
timestamp 1663859327
transform 1 0 40768 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_384
timestamp 1663859327
transform 1 0 44352 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_48_388
timestamp 1663859327
transform 1 0 44800 0 1 40768
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_48_392
timestamp 1663859327
transform 1 0 45248 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_48_408
timestamp 1663859327
transform 1 0 47040 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_48_416
timestamp 1663859327
transform 1 0 47936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_2
timestamp 1663859327
transform 1 0 1568 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_8
timestamp 1663859327
transform 1 0 2240 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_12
timestamp 1663859327
transform 1 0 2688 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_16
timestamp 1663859327
transform 1 0 3136 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_20
timestamp 1663859327
transform 1 0 3584 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_24
timestamp 1663859327
transform 1 0 4032 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_28
timestamp 1663859327
transform 1 0 4480 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_32
timestamp 1663859327
transform 1 0 4928 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_36
timestamp 1663859327
transform 1 0 5376 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_40
timestamp 1663859327
transform 1 0 5824 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_44
timestamp 1663859327
transform 1 0 6272 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_52
timestamp 1663859327
transform 1 0 7168 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_60
timestamp 1663859327
transform 1 0 8064 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_70
timestamp 1663859327
transform 1 0 9184 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_73
timestamp 1663859327
transform 1 0 9520 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_79
timestamp 1663859327
transform 1 0 10192 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_110
timestamp 1663859327
transform 1 0 13664 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_141
timestamp 1663859327
transform 1 0 17136 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_144
timestamp 1663859327
transform 1 0 17472 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_155
timestamp 1663859327
transform 1 0 18704 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_188
timestamp 1663859327
transform 1 0 22400 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_209
timestamp 1663859327
transform 1 0 24752 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_215
timestamp 1663859327
transform 1 0 25424 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_245
timestamp 1663859327
transform 1 0 28784 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_270
timestamp 1663859327
transform 1 0 31584 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_282
timestamp 1663859327
transform 1 0 32928 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_286
timestamp 1663859327
transform 1 0 33376 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_295
timestamp 1663859327
transform 1 0 34384 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_303
timestamp 1663859327
transform 1 0 35280 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_307
timestamp 1663859327
transform 1 0 35728 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_311
timestamp 1663859327
transform 1 0 36176 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_315
timestamp 1663859327
transform 1 0 36624 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_319
timestamp 1663859327
transform 1 0 37072 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_323
timestamp 1663859327
transform 1 0 37520 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_327
timestamp 1663859327
transform 1 0 37968 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_331
timestamp 1663859327
transform 1 0 38416 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_335
timestamp 1663859327
transform 1 0 38864 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_339
timestamp 1663859327
transform 1 0 39312 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_343
timestamp 1663859327
transform 1 0 39760 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_49_347
timestamp 1663859327
transform 1 0 40208 0 -1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_351
timestamp 1663859327
transform 1 0 40656 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_49_357
timestamp 1663859327
transform 1 0 41328 0 -1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_49_360
timestamp 1663859327
transform 1 0 41664 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_49_392
timestamp 1663859327
transform 1 0 45248 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_49_408
timestamp 1663859327
transform 1 0 47040 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_49_416
timestamp 1663859327
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_2
timestamp 1663859327
transform 1 0 1568 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_7
timestamp 1663859327
transform 1 0 2128 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_11
timestamp 1663859327
transform 1 0 2576 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_14
timestamp 1663859327
transform 1 0 2912 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_18
timestamp 1663859327
transform 1 0 3360 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_22
timestamp 1663859327
transform 1 0 3808 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_26
timestamp 1663859327
transform 1 0 4256 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_30
timestamp 1663859327
transform 1 0 4704 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_34
timestamp 1663859327
transform 1 0 5152 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_37
timestamp 1663859327
transform 1 0 5488 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_39
timestamp 1663859327
transform 1 0 5712 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_42
timestamp 1663859327
transform 1 0 6048 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_46
timestamp 1663859327
transform 1 0 6496 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_50
timestamp 1663859327
transform 1 0 6944 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_54
timestamp 1663859327
transform 1 0 7392 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_58
timestamp 1663859327
transform 1 0 7840 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_66
timestamp 1663859327
transform 1 0 8736 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_74
timestamp 1663859327
transform 1 0 9632 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_105
timestamp 1663859327
transform 1 0 13104 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_108
timestamp 1663859327
transform 1 0 13440 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_114
timestamp 1663859327
transform 1 0 14112 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_145
timestamp 1663859327
transform 1 0 17584 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_176
timestamp 1663859327
transform 1 0 21056 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_179
timestamp 1663859327
transform 1 0 21392 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_209
timestamp 1663859327
transform 1 0 24752 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_240
timestamp 1663859327
transform 1 0 28224 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_247
timestamp 1663859327
transform 1 0 29008 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_250
timestamp 1663859327
transform 1 0 29344 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_263
timestamp 1663859327
transform 1 0 30800 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_275
timestamp 1663859327
transform 1 0 32144 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_285
timestamp 1663859327
transform 1 0 33264 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_293
timestamp 1663859327
transform 1 0 34160 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_297
timestamp 1663859327
transform 1 0 34608 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_301
timestamp 1663859327
transform 1 0 35056 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_305
timestamp 1663859327
transform 1 0 35504 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_309
timestamp 1663859327
transform 1 0 35952 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_313
timestamp 1663859327
transform 1 0 36400 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_317
timestamp 1663859327
transform 1 0 36848 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_50_321
timestamp 1663859327
transform 1 0 37296 0 1 42336
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_324
timestamp 1663859327
transform 1 0 37632 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_328
timestamp 1663859327
transform 1 0 38080 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_332
timestamp 1663859327
transform 1 0 38528 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_336
timestamp 1663859327
transform 1 0 38976 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_340
timestamp 1663859327
transform 1 0 39424 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_344
timestamp 1663859327
transform 1 0 39872 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_348
timestamp 1663859327
transform 1 0 40320 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_50_352
timestamp 1663859327
transform 1 0 40768 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_384
timestamp 1663859327
transform 1 0 44352 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_50_388
timestamp 1663859327
transform 1 0 44800 0 1 42336
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_50_392
timestamp 1663859327
transform 1 0 45248 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_50_408
timestamp 1663859327
transform 1 0 47040 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_50_416
timestamp 1663859327
transform 1 0 47936 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_2
timestamp 1663859327
transform 1 0 1568 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_6
timestamp 1663859327
transform 1 0 2016 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_10
timestamp 1663859327
transform 1 0 2464 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_14
timestamp 1663859327
transform 1 0 2912 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_18
timestamp 1663859327
transform 1 0 3360 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_22
timestamp 1663859327
transform 1 0 3808 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_26
timestamp 1663859327
transform 1 0 4256 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_30
timestamp 1663859327
transform 1 0 4704 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_34
timestamp 1663859327
transform 1 0 5152 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_38
timestamp 1663859327
transform 1 0 5600 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_42
timestamp 1663859327
transform 1 0 6048 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_46
timestamp 1663859327
transform 1 0 6496 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_50
timestamp 1663859327
transform 1 0 6944 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_54
timestamp 1663859327
transform 1 0 7392 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_58
timestamp 1663859327
transform 1 0 7840 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_62
timestamp 1663859327
transform 1 0 8288 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_66
timestamp 1663859327
transform 1 0 8736 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_70
timestamp 1663859327
transform 1 0 9184 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_73
timestamp 1663859327
transform 1 0 9520 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_77
timestamp 1663859327
transform 1 0 9968 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_85
timestamp 1663859327
transform 1 0 10864 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_95
timestamp 1663859327
transform 1 0 11984 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_110
timestamp 1663859327
transform 1 0 13664 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_141
timestamp 1663859327
transform 1 0 17136 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_144
timestamp 1663859327
transform 1 0 17472 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_160
timestamp 1663859327
transform 1 0 19264 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_191
timestamp 1663859327
transform 1 0 22736 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_211
timestamp 1663859327
transform 1 0 24976 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_215
timestamp 1663859327
transform 1 0 25424 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_245
timestamp 1663859327
transform 1 0 28784 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_258
timestamp 1663859327
transform 1 0 30240 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_269
timestamp 1663859327
transform 1 0 31472 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_278
timestamp 1663859327
transform 1 0 32480 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_282
timestamp 1663859327
transform 1 0 32928 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_286
timestamp 1663859327
transform 1 0 33376 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_289
timestamp 1663859327
transform 1 0 33712 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_293
timestamp 1663859327
transform 1 0 34160 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_297
timestamp 1663859327
transform 1 0 34608 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_301
timestamp 1663859327
transform 1 0 35056 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_305
timestamp 1663859327
transform 1 0 35504 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_309
timestamp 1663859327
transform 1 0 35952 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_313
timestamp 1663859327
transform 1 0 36400 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_317
timestamp 1663859327
transform 1 0 36848 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_321
timestamp 1663859327
transform 1 0 37296 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_325
timestamp 1663859327
transform 1 0 37744 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_329
timestamp 1663859327
transform 1 0 38192 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_333
timestamp 1663859327
transform 1 0 38640 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_337
timestamp 1663859327
transform 1 0 39088 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_341
timestamp 1663859327
transform 1 0 39536 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_345
timestamp 1663859327
transform 1 0 39984 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_349
timestamp 1663859327
transform 1 0 40432 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_353
timestamp 1663859327
transform 1 0 40880 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_51_357
timestamp 1663859327
transform 1 0 41328 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_51_389
timestamp 1663859327
transform 1 0 44912 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_51_405
timestamp 1663859327
transform 1 0 46704 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_51_411
timestamp 1663859327
transform 1 0 47376 0 -1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_51_419
timestamp 1663859327
transform 1 0 48272 0 -1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_2
timestamp 1663859327
transform 1 0 1568 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_17
timestamp 1663859327
transform 1 0 3248 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_19
timestamp 1663859327
transform 1 0 3472 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_22
timestamp 1663859327
transform 1 0 3808 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_26
timestamp 1663859327
transform 1 0 4256 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_30
timestamp 1663859327
transform 1 0 4704 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_34
timestamp 1663859327
transform 1 0 5152 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_37
timestamp 1663859327
transform 1 0 5488 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_41
timestamp 1663859327
transform 1 0 5936 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_45
timestamp 1663859327
transform 1 0 6384 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_49
timestamp 1663859327
transform 1 0 6832 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_53
timestamp 1663859327
transform 1 0 7280 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_57
timestamp 1663859327
transform 1 0 7728 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_61
timestamp 1663859327
transform 1 0 8176 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_65
timestamp 1663859327
transform 1 0 8624 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_69
timestamp 1663859327
transform 1 0 9072 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_73
timestamp 1663859327
transform 1 0 9520 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_77
timestamp 1663859327
transform 1 0 9968 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_85
timestamp 1663859327
transform 1 0 10864 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_95
timestamp 1663859327
transform 1 0 11984 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_105
timestamp 1663859327
transform 1 0 13104 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_108
timestamp 1663859327
transform 1 0 13440 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_114
timestamp 1663859327
transform 1 0 14112 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_145
timestamp 1663859327
transform 1 0 17584 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_176
timestamp 1663859327
transform 1 0 21056 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_179
timestamp 1663859327
transform 1 0 21392 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_209
timestamp 1663859327
transform 1 0 24752 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_240
timestamp 1663859327
transform 1 0 28224 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_247
timestamp 1663859327
transform 1 0 29008 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_250
timestamp 1663859327
transform 1 0 29344 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_259
timestamp 1663859327
transform 1 0 30352 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_269
timestamp 1663859327
transform 1 0 31472 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_277
timestamp 1663859327
transform 1 0 32368 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_281
timestamp 1663859327
transform 1 0 32816 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_285
timestamp 1663859327
transform 1 0 33264 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_289
timestamp 1663859327
transform 1 0 33712 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_293
timestamp 1663859327
transform 1 0 34160 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_297
timestamp 1663859327
transform 1 0 34608 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_301
timestamp 1663859327
transform 1 0 35056 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_305
timestamp 1663859327
transform 1 0 35504 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_309
timestamp 1663859327
transform 1 0 35952 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_313
timestamp 1663859327
transform 1 0 36400 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_317
timestamp 1663859327
transform 1 0 36848 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_52_321
timestamp 1663859327
transform 1 0 37296 0 1 43904
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_324
timestamp 1663859327
transform 1 0 37632 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_328
timestamp 1663859327
transform 1 0 38080 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_332
timestamp 1663859327
transform 1 0 38528 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_336
timestamp 1663859327
transform 1 0 38976 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_340
timestamp 1663859327
transform 1 0 39424 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_344
timestamp 1663859327
transform 1 0 39872 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_52_348
timestamp 1663859327
transform 1 0 40320 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_380
timestamp 1663859327
transform 1 0 43904 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_52_388
timestamp 1663859327
transform 1 0 44800 0 1 43904
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_52_392
timestamp 1663859327
transform 1 0 45248 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_52_408
timestamp 1663859327
transform 1 0 47040 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_52_416
timestamp 1663859327
transform 1 0 47936 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_2
timestamp 1663859327
transform 1 0 1568 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_7
timestamp 1663859327
transform 1 0 2128 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_13
timestamp 1663859327
transform 1 0 2800 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_19
timestamp 1663859327
transform 1 0 3472 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_23
timestamp 1663859327
transform 1 0 3920 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_26
timestamp 1663859327
transform 1 0 4256 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_30
timestamp 1663859327
transform 1 0 4704 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_34
timestamp 1663859327
transform 1 0 5152 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_38
timestamp 1663859327
transform 1 0 5600 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_42
timestamp 1663859327
transform 1 0 6048 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_46
timestamp 1663859327
transform 1 0 6496 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_50
timestamp 1663859327
transform 1 0 6944 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_54
timestamp 1663859327
transform 1 0 7392 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_58
timestamp 1663859327
transform 1 0 7840 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_62
timestamp 1663859327
transform 1 0 8288 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_66
timestamp 1663859327
transform 1 0 8736 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_70
timestamp 1663859327
transform 1 0 9184 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_73
timestamp 1663859327
transform 1 0 9520 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_76
timestamp 1663859327
transform 1 0 9856 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_80
timestamp 1663859327
transform 1 0 10304 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_84
timestamp 1663859327
transform 1 0 10752 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_92
timestamp 1663859327
transform 1 0 11648 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_100
timestamp 1663859327
transform 1 0 12544 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_110
timestamp 1663859327
transform 1 0 13664 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_141
timestamp 1663859327
transform 1 0 17136 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_144
timestamp 1663859327
transform 1 0 17472 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_159
timestamp 1663859327
transform 1 0 19152 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_190
timestamp 1663859327
transform 1 0 22624 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_208
timestamp 1663859327
transform 1 0 24640 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_212
timestamp 1663859327
transform 1 0 25088 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_215
timestamp 1663859327
transform 1 0 25424 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_231
timestamp 1663859327
transform 1 0 27216 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_243
timestamp 1663859327
transform 1 0 28560 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_253
timestamp 1663859327
transform 1 0 29680 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_261
timestamp 1663859327
transform 1 0 30576 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_267
timestamp 1663859327
transform 1 0 31248 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_271
timestamp 1663859327
transform 1 0 31696 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_275
timestamp 1663859327
transform 1 0 32144 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_279
timestamp 1663859327
transform 1 0 32592 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_283
timestamp 1663859327
transform 1 0 33040 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_286
timestamp 1663859327
transform 1 0 33376 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_289
timestamp 1663859327
transform 1 0 33712 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_293
timestamp 1663859327
transform 1 0 34160 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_297
timestamp 1663859327
transform 1 0 34608 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_301
timestamp 1663859327
transform 1 0 35056 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_305
timestamp 1663859327
transform 1 0 35504 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_309
timestamp 1663859327
transform 1 0 35952 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_313
timestamp 1663859327
transform 1 0 36400 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_317
timestamp 1663859327
transform 1 0 36848 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_321
timestamp 1663859327
transform 1 0 37296 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_325
timestamp 1663859327
transform 1 0 37744 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_329
timestamp 1663859327
transform 1 0 38192 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_333
timestamp 1663859327
transform 1 0 38640 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_337
timestamp 1663859327
transform 1 0 39088 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_341
timestamp 1663859327
transform 1 0 39536 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_345
timestamp 1663859327
transform 1 0 39984 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_349
timestamp 1663859327
transform 1 0 40432 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_353
timestamp 1663859327
transform 1 0 40880 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_53_357
timestamp 1663859327
transform 1 0 41328 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_53_389
timestamp 1663859327
transform 1 0 44912 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_53_405
timestamp 1663859327
transform 1 0 46704 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_53_413
timestamp 1663859327
transform 1 0 47600 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_53_417
timestamp 1663859327
transform 1 0 48048 0 -1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_53_419
timestamp 1663859327
transform 1 0 48272 0 -1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_2
timestamp 1663859327
transform 1 0 1568 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_9
timestamp 1663859327
transform 1 0 2352 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_15
timestamp 1663859327
transform 1 0 3024 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_19
timestamp 1663859327
transform 1 0 3472 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_34
timestamp 1663859327
transform 1 0 5152 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_37
timestamp 1663859327
transform 1 0 5488 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_41
timestamp 1663859327
transform 1 0 5936 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_45
timestamp 1663859327
transform 1 0 6384 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_49
timestamp 1663859327
transform 1 0 6832 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_53
timestamp 1663859327
transform 1 0 7280 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_59
timestamp 1663859327
transform 1 0 7952 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_63
timestamp 1663859327
transform 1 0 8400 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_69
timestamp 1663859327
transform 1 0 9072 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_72
timestamp 1663859327
transform 1 0 9408 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_76
timestamp 1663859327
transform 1 0 9856 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_82
timestamp 1663859327
transform 1 0 10528 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_88
timestamp 1663859327
transform 1 0 11200 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_96
timestamp 1663859327
transform 1 0 12096 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_104
timestamp 1663859327
transform 1 0 12992 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_107
timestamp 1663859327
transform 1 0 13328 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_134
timestamp 1663859327
transform 1 0 16352 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_136
timestamp 1663859327
transform 1 0 16576 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_139
timestamp 1663859327
transform 1 0 16912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_142
timestamp 1663859327
transform 1 0 17248 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_144
timestamp 1663859327
transform 1 0 17472 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_174
timestamp 1663859327
transform 1 0 20832 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_177
timestamp 1663859327
transform 1 0 21168 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_207
timestamp 1663859327
transform 1 0 24528 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_209
timestamp 1663859327
transform 1 0 24752 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_212
timestamp 1663859327
transform 1 0 25088 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_226
timestamp 1663859327
transform 1 0 26656 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_238
timestamp 1663859327
transform 1 0 28000 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_244
timestamp 1663859327
transform 1 0 28672 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_247
timestamp 1663859327
transform 1 0 29008 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_254
timestamp 1663859327
transform 1 0 29792 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_260
timestamp 1663859327
transform 1 0 30464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_264
timestamp 1663859327
transform 1 0 30912 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_271
timestamp 1663859327
transform 1 0 31696 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_277
timestamp 1663859327
transform 1 0 32368 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_279
timestamp 1663859327
transform 1 0 32592 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_282
timestamp 1663859327
transform 1 0 32928 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_297
timestamp 1663859327
transform 1 0 34608 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_299
timestamp 1663859327
transform 1 0 34832 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_314
timestamp 1663859327
transform 1 0 36512 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_317
timestamp 1663859327
transform 1 0 36848 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_320
timestamp 1663859327
transform 1 0 37184 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_324
timestamp 1663859327
transform 1 0 37632 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_329
timestamp 1663859327
transform 1 0 38192 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_333
timestamp 1663859327
transform 1 0 38640 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_337
timestamp 1663859327
transform 1 0 39088 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_341
timestamp 1663859327
transform 1 0 39536 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_347
timestamp 1663859327
transform 1 0 40208 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_349
timestamp 1663859327
transform 1 0 40432 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_352
timestamp 1663859327
transform 1 0 40768 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_355
timestamp 1663859327
transform 1 0 41104 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_359
timestamp 1663859327
transform 1 0 41552 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_363
timestamp 1663859327
transform 1 0 42000 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_54_371
timestamp 1663859327
transform 1 0 42896 0 1 45472
box 0 -60 224 844
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_377
timestamp 1663859327
transform 1 0 43568 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_54_387
timestamp 1663859327
transform 1 0 44688 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_54_403
timestamp 1663859327
transform 1 0 46480 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_54_411
timestamp 1663859327
transform 1 0 47376 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_54_419
timestamp 1663859327
transform 1 0 48272 0 1 45472
box 0 -60 112 844
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_0 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_1
timestamp 1663859327
transform -1 0 48608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_2
timestamp 1663859327
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_3
timestamp 1663859327
transform -1 0 48608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_4
timestamp 1663859327
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_5
timestamp 1663859327
transform -1 0 48608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_6
timestamp 1663859327
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_7
timestamp 1663859327
transform -1 0 48608 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_8
timestamp 1663859327
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_9
timestamp 1663859327
transform -1 0 48608 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_10
timestamp 1663859327
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_11
timestamp 1663859327
transform -1 0 48608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_12
timestamp 1663859327
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_13
timestamp 1663859327
transform -1 0 48608 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_14
timestamp 1663859327
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_15
timestamp 1663859327
transform -1 0 48608 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_16
timestamp 1663859327
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_17
timestamp 1663859327
transform -1 0 48608 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_18
timestamp 1663859327
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_19
timestamp 1663859327
transform -1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_20
timestamp 1663859327
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_21
timestamp 1663859327
transform -1 0 48608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_22
timestamp 1663859327
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_23
timestamp 1663859327
transform -1 0 48608 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_24
timestamp 1663859327
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_25
timestamp 1663859327
transform -1 0 48608 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_26
timestamp 1663859327
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_27
timestamp 1663859327
transform -1 0 48608 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_28
timestamp 1663859327
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_29
timestamp 1663859327
transform -1 0 48608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_30
timestamp 1663859327
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_31
timestamp 1663859327
transform -1 0 48608 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_32
timestamp 1663859327
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_33
timestamp 1663859327
transform -1 0 48608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_34
timestamp 1663859327
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_35
timestamp 1663859327
transform -1 0 48608 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_36
timestamp 1663859327
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_37
timestamp 1663859327
transform -1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_38
timestamp 1663859327
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_39
timestamp 1663859327
transform -1 0 48608 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_40
timestamp 1663859327
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_41
timestamp 1663859327
transform -1 0 48608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_42
timestamp 1663859327
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_43
timestamp 1663859327
transform -1 0 48608 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_44
timestamp 1663859327
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_45
timestamp 1663859327
transform -1 0 48608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_46
timestamp 1663859327
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_47
timestamp 1663859327
transform -1 0 48608 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_48
timestamp 1663859327
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_49
timestamp 1663859327
transform -1 0 48608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_50
timestamp 1663859327
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_51
timestamp 1663859327
transform -1 0 48608 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_52
timestamp 1663859327
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_53
timestamp 1663859327
transform -1 0 48608 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_54
timestamp 1663859327
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_55
timestamp 1663859327
transform -1 0 48608 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_56
timestamp 1663859327
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_57
timestamp 1663859327
transform -1 0 48608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_58
timestamp 1663859327
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_59
timestamp 1663859327
transform -1 0 48608 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_60
timestamp 1663859327
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_61
timestamp 1663859327
transform -1 0 48608 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_62
timestamp 1663859327
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_63
timestamp 1663859327
transform -1 0 48608 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_64
timestamp 1663859327
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_65
timestamp 1663859327
transform -1 0 48608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_66
timestamp 1663859327
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_67
timestamp 1663859327
transform -1 0 48608 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_68
timestamp 1663859327
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_69
timestamp 1663859327
transform -1 0 48608 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_70
timestamp 1663859327
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_71
timestamp 1663859327
transform -1 0 48608 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_72
timestamp 1663859327
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_73
timestamp 1663859327
transform -1 0 48608 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_74
timestamp 1663859327
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_75
timestamp 1663859327
transform -1 0 48608 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_76
timestamp 1663859327
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_77
timestamp 1663859327
transform -1 0 48608 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_78
timestamp 1663859327
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_79
timestamp 1663859327
transform -1 0 48608 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_80
timestamp 1663859327
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_81
timestamp 1663859327
transform -1 0 48608 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_82
timestamp 1663859327
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_83
timestamp 1663859327
transform -1 0 48608 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_84
timestamp 1663859327
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_85
timestamp 1663859327
transform -1 0 48608 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_86
timestamp 1663859327
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_87
timestamp 1663859327
transform -1 0 48608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_88
timestamp 1663859327
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_89
timestamp 1663859327
transform -1 0 48608 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_90
timestamp 1663859327
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_91
timestamp 1663859327
transform -1 0 48608 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_92
timestamp 1663859327
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_93
timestamp 1663859327
transform -1 0 48608 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_94
timestamp 1663859327
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_95
timestamp 1663859327
transform -1 0 48608 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_96
timestamp 1663859327
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_97
timestamp 1663859327
transform -1 0 48608 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_98
timestamp 1663859327
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_99
timestamp 1663859327
transform -1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_100
timestamp 1663859327
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_101
timestamp 1663859327
transform -1 0 48608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_102
timestamp 1663859327
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_103
timestamp 1663859327
transform -1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_104
timestamp 1663859327
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_105
timestamp 1663859327
transform -1 0 48608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_106
timestamp 1663859327
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_107
timestamp 1663859327
transform -1 0 48608 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_108
timestamp 1663859327
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_109
timestamp 1663859327
transform -1 0 48608 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_110 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 5264 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_111
timestamp 1663859327
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_112
timestamp 1663859327
transform 1 0 13104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_113
timestamp 1663859327
transform 1 0 17024 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_114
timestamp 1663859327
transform 1 0 20944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_115
timestamp 1663859327
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_116
timestamp 1663859327
transform 1 0 28784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_117
timestamp 1663859327
transform 1 0 32704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_118
timestamp 1663859327
transform 1 0 36624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_119
timestamp 1663859327
transform 1 0 40544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_120
timestamp 1663859327
transform 1 0 44464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_121
timestamp 1663859327
transform 1 0 9296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_122
timestamp 1663859327
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_123
timestamp 1663859327
transform 1 0 25200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_124
timestamp 1663859327
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_125
timestamp 1663859327
transform 1 0 41104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_126
timestamp 1663859327
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_127
timestamp 1663859327
transform 1 0 13216 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_128
timestamp 1663859327
transform 1 0 21168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_129
timestamp 1663859327
transform 1 0 29120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_130
timestamp 1663859327
transform 1 0 37072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_131
timestamp 1663859327
transform 1 0 45024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_132
timestamp 1663859327
transform 1 0 9296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_133
timestamp 1663859327
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_134
timestamp 1663859327
transform 1 0 25200 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_135
timestamp 1663859327
transform 1 0 33152 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_136
timestamp 1663859327
transform 1 0 41104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_137
timestamp 1663859327
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_138
timestamp 1663859327
transform 1 0 13216 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_139
timestamp 1663859327
transform 1 0 21168 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_140
timestamp 1663859327
transform 1 0 29120 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_141
timestamp 1663859327
transform 1 0 37072 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_142
timestamp 1663859327
transform 1 0 45024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_143
timestamp 1663859327
transform 1 0 9296 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_144
timestamp 1663859327
transform 1 0 17248 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_145
timestamp 1663859327
transform 1 0 25200 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_146
timestamp 1663859327
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_147
timestamp 1663859327
transform 1 0 41104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_148
timestamp 1663859327
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_149
timestamp 1663859327
transform 1 0 13216 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_150
timestamp 1663859327
transform 1 0 21168 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_151
timestamp 1663859327
transform 1 0 29120 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_152
timestamp 1663859327
transform 1 0 37072 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_153
timestamp 1663859327
transform 1 0 45024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_154
timestamp 1663859327
transform 1 0 9296 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_155
timestamp 1663859327
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_156
timestamp 1663859327
transform 1 0 25200 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_157
timestamp 1663859327
transform 1 0 33152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_158
timestamp 1663859327
transform 1 0 41104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_159
timestamp 1663859327
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_160
timestamp 1663859327
transform 1 0 13216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_161
timestamp 1663859327
transform 1 0 21168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_162
timestamp 1663859327
transform 1 0 29120 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_163
timestamp 1663859327
transform 1 0 37072 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_164
timestamp 1663859327
transform 1 0 45024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_165
timestamp 1663859327
transform 1 0 9296 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_166
timestamp 1663859327
transform 1 0 17248 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_167
timestamp 1663859327
transform 1 0 25200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_168
timestamp 1663859327
transform 1 0 33152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_169
timestamp 1663859327
transform 1 0 41104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_170
timestamp 1663859327
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_171
timestamp 1663859327
transform 1 0 13216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_172
timestamp 1663859327
transform 1 0 21168 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_173
timestamp 1663859327
transform 1 0 29120 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_174
timestamp 1663859327
transform 1 0 37072 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_175
timestamp 1663859327
transform 1 0 45024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_176
timestamp 1663859327
transform 1 0 9296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_177
timestamp 1663859327
transform 1 0 17248 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_178
timestamp 1663859327
transform 1 0 25200 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_179
timestamp 1663859327
transform 1 0 33152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_180
timestamp 1663859327
transform 1 0 41104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_181
timestamp 1663859327
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_182
timestamp 1663859327
transform 1 0 13216 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_183
timestamp 1663859327
transform 1 0 21168 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_184
timestamp 1663859327
transform 1 0 29120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_185
timestamp 1663859327
transform 1 0 37072 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_186
timestamp 1663859327
transform 1 0 45024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_187
timestamp 1663859327
transform 1 0 9296 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_188
timestamp 1663859327
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_189
timestamp 1663859327
transform 1 0 25200 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_190
timestamp 1663859327
transform 1 0 33152 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_191
timestamp 1663859327
transform 1 0 41104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_192
timestamp 1663859327
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_193
timestamp 1663859327
transform 1 0 13216 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_194
timestamp 1663859327
transform 1 0 21168 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_195
timestamp 1663859327
transform 1 0 29120 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_196
timestamp 1663859327
transform 1 0 37072 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_197
timestamp 1663859327
transform 1 0 45024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_198
timestamp 1663859327
transform 1 0 9296 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_199
timestamp 1663859327
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_200
timestamp 1663859327
transform 1 0 25200 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_201
timestamp 1663859327
transform 1 0 33152 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_202
timestamp 1663859327
transform 1 0 41104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_203
timestamp 1663859327
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_204
timestamp 1663859327
transform 1 0 13216 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_205
timestamp 1663859327
transform 1 0 21168 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_206
timestamp 1663859327
transform 1 0 29120 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_207
timestamp 1663859327
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_208
timestamp 1663859327
transform 1 0 45024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_209
timestamp 1663859327
transform 1 0 9296 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_210
timestamp 1663859327
transform 1 0 17248 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_211
timestamp 1663859327
transform 1 0 25200 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_212
timestamp 1663859327
transform 1 0 33152 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_213
timestamp 1663859327
transform 1 0 41104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_214
timestamp 1663859327
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_215
timestamp 1663859327
transform 1 0 13216 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_216
timestamp 1663859327
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_217
timestamp 1663859327
transform 1 0 29120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_218
timestamp 1663859327
transform 1 0 37072 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_219
timestamp 1663859327
transform 1 0 45024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_220
timestamp 1663859327
transform 1 0 9296 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_221
timestamp 1663859327
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_222
timestamp 1663859327
transform 1 0 25200 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_223
timestamp 1663859327
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_224
timestamp 1663859327
transform 1 0 41104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_225
timestamp 1663859327
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_226
timestamp 1663859327
transform 1 0 13216 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_227
timestamp 1663859327
transform 1 0 21168 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_228
timestamp 1663859327
transform 1 0 29120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_229
timestamp 1663859327
transform 1 0 37072 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_230
timestamp 1663859327
transform 1 0 45024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_231
timestamp 1663859327
transform 1 0 9296 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_232
timestamp 1663859327
transform 1 0 17248 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_233
timestamp 1663859327
transform 1 0 25200 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_234
timestamp 1663859327
transform 1 0 33152 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_235
timestamp 1663859327
transform 1 0 41104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_236
timestamp 1663859327
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_237
timestamp 1663859327
transform 1 0 13216 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_238
timestamp 1663859327
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_239
timestamp 1663859327
transform 1 0 29120 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_240
timestamp 1663859327
transform 1 0 37072 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_241
timestamp 1663859327
transform 1 0 45024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_242
timestamp 1663859327
transform 1 0 9296 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_243
timestamp 1663859327
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_244
timestamp 1663859327
transform 1 0 25200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_245
timestamp 1663859327
transform 1 0 33152 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_246
timestamp 1663859327
transform 1 0 41104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_247
timestamp 1663859327
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_248
timestamp 1663859327
transform 1 0 13216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_249
timestamp 1663859327
transform 1 0 21168 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_250
timestamp 1663859327
transform 1 0 29120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_251
timestamp 1663859327
transform 1 0 37072 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_252
timestamp 1663859327
transform 1 0 45024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_253
timestamp 1663859327
transform 1 0 9296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_254
timestamp 1663859327
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_255
timestamp 1663859327
transform 1 0 25200 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_256
timestamp 1663859327
transform 1 0 33152 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_257
timestamp 1663859327
transform 1 0 41104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_258
timestamp 1663859327
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_259
timestamp 1663859327
transform 1 0 13216 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_260
timestamp 1663859327
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_261
timestamp 1663859327
transform 1 0 29120 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_262
timestamp 1663859327
transform 1 0 37072 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_263
timestamp 1663859327
transform 1 0 45024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_264
timestamp 1663859327
transform 1 0 9296 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_265
timestamp 1663859327
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_266
timestamp 1663859327
transform 1 0 25200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_267
timestamp 1663859327
transform 1 0 33152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_268
timestamp 1663859327
transform 1 0 41104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_269
timestamp 1663859327
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_270
timestamp 1663859327
transform 1 0 13216 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_271
timestamp 1663859327
transform 1 0 21168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_272
timestamp 1663859327
transform 1 0 29120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_273
timestamp 1663859327
transform 1 0 37072 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_274
timestamp 1663859327
transform 1 0 45024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_275
timestamp 1663859327
transform 1 0 9296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_276
timestamp 1663859327
transform 1 0 17248 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_277
timestamp 1663859327
transform 1 0 25200 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_278
timestamp 1663859327
transform 1 0 33152 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_279
timestamp 1663859327
transform 1 0 41104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_280
timestamp 1663859327
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_281
timestamp 1663859327
transform 1 0 13216 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_282
timestamp 1663859327
transform 1 0 21168 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_283
timestamp 1663859327
transform 1 0 29120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_284
timestamp 1663859327
transform 1 0 37072 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_285
timestamp 1663859327
transform 1 0 45024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_286
timestamp 1663859327
transform 1 0 9296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_287
timestamp 1663859327
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_288
timestamp 1663859327
transform 1 0 25200 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_289
timestamp 1663859327
transform 1 0 33152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_290
timestamp 1663859327
transform 1 0 41104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_291
timestamp 1663859327
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_292
timestamp 1663859327
transform 1 0 13216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_293
timestamp 1663859327
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_294
timestamp 1663859327
transform 1 0 29120 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_295
timestamp 1663859327
transform 1 0 37072 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_296
timestamp 1663859327
transform 1 0 45024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_297
timestamp 1663859327
transform 1 0 9296 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_298
timestamp 1663859327
transform 1 0 17248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_299
timestamp 1663859327
transform 1 0 25200 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_300
timestamp 1663859327
transform 1 0 33152 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_301
timestamp 1663859327
transform 1 0 41104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_302
timestamp 1663859327
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_303
timestamp 1663859327
transform 1 0 13216 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_304
timestamp 1663859327
transform 1 0 21168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_305
timestamp 1663859327
transform 1 0 29120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_306
timestamp 1663859327
transform 1 0 37072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_307
timestamp 1663859327
transform 1 0 45024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_308
timestamp 1663859327
transform 1 0 9296 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_309
timestamp 1663859327
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_310
timestamp 1663859327
transform 1 0 25200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_311
timestamp 1663859327
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_312
timestamp 1663859327
transform 1 0 41104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_313
timestamp 1663859327
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_314
timestamp 1663859327
transform 1 0 13216 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_315
timestamp 1663859327
transform 1 0 21168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_316
timestamp 1663859327
transform 1 0 29120 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_317
timestamp 1663859327
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_318
timestamp 1663859327
transform 1 0 45024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_319
timestamp 1663859327
transform 1 0 9296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_320
timestamp 1663859327
transform 1 0 17248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_321
timestamp 1663859327
transform 1 0 25200 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_322
timestamp 1663859327
transform 1 0 33152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_323
timestamp 1663859327
transform 1 0 41104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_324
timestamp 1663859327
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_325
timestamp 1663859327
transform 1 0 13216 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_326
timestamp 1663859327
transform 1 0 21168 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_327
timestamp 1663859327
transform 1 0 29120 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_328
timestamp 1663859327
transform 1 0 37072 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_329
timestamp 1663859327
transform 1 0 45024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_330
timestamp 1663859327
transform 1 0 9296 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_331
timestamp 1663859327
transform 1 0 17248 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_332
timestamp 1663859327
transform 1 0 25200 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_333
timestamp 1663859327
transform 1 0 33152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_334
timestamp 1663859327
transform 1 0 41104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_335
timestamp 1663859327
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_336
timestamp 1663859327
transform 1 0 13216 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_337
timestamp 1663859327
transform 1 0 21168 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_338
timestamp 1663859327
transform 1 0 29120 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_339
timestamp 1663859327
transform 1 0 37072 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_340
timestamp 1663859327
transform 1 0 45024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_341
timestamp 1663859327
transform 1 0 9296 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_342
timestamp 1663859327
transform 1 0 17248 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_343
timestamp 1663859327
transform 1 0 25200 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_344
timestamp 1663859327
transform 1 0 33152 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_345
timestamp 1663859327
transform 1 0 41104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_346
timestamp 1663859327
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_347
timestamp 1663859327
transform 1 0 13216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_348
timestamp 1663859327
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_349
timestamp 1663859327
transform 1 0 29120 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_350
timestamp 1663859327
transform 1 0 37072 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_351
timestamp 1663859327
transform 1 0 45024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_352
timestamp 1663859327
transform 1 0 9296 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_353
timestamp 1663859327
transform 1 0 17248 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_354
timestamp 1663859327
transform 1 0 25200 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_355
timestamp 1663859327
transform 1 0 33152 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_356
timestamp 1663859327
transform 1 0 41104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_357
timestamp 1663859327
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_358
timestamp 1663859327
transform 1 0 13216 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_359
timestamp 1663859327
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_360
timestamp 1663859327
transform 1 0 29120 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_361
timestamp 1663859327
transform 1 0 37072 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_362
timestamp 1663859327
transform 1 0 45024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_363
timestamp 1663859327
transform 1 0 9296 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_364
timestamp 1663859327
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_365
timestamp 1663859327
transform 1 0 25200 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_366
timestamp 1663859327
transform 1 0 33152 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_367
timestamp 1663859327
transform 1 0 41104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_368
timestamp 1663859327
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_369
timestamp 1663859327
transform 1 0 13216 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_370
timestamp 1663859327
transform 1 0 21168 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_371
timestamp 1663859327
transform 1 0 29120 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_372
timestamp 1663859327
transform 1 0 37072 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_373
timestamp 1663859327
transform 1 0 45024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_374
timestamp 1663859327
transform 1 0 9296 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_375
timestamp 1663859327
transform 1 0 17248 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_376
timestamp 1663859327
transform 1 0 25200 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_377
timestamp 1663859327
transform 1 0 33152 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_378
timestamp 1663859327
transform 1 0 41104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_379
timestamp 1663859327
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_380
timestamp 1663859327
transform 1 0 13216 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_381
timestamp 1663859327
transform 1 0 21168 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_382
timestamp 1663859327
transform 1 0 29120 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_383
timestamp 1663859327
transform 1 0 37072 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_384
timestamp 1663859327
transform 1 0 45024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_385
timestamp 1663859327
transform 1 0 9296 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_386
timestamp 1663859327
transform 1 0 17248 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_387
timestamp 1663859327
transform 1 0 25200 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_388
timestamp 1663859327
transform 1 0 33152 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_389
timestamp 1663859327
transform 1 0 41104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_390
timestamp 1663859327
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_391
timestamp 1663859327
transform 1 0 13216 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_392
timestamp 1663859327
transform 1 0 21168 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_393
timestamp 1663859327
transform 1 0 29120 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_394
timestamp 1663859327
transform 1 0 37072 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_395
timestamp 1663859327
transform 1 0 45024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_396
timestamp 1663859327
transform 1 0 9296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_397
timestamp 1663859327
transform 1 0 17248 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_398
timestamp 1663859327
transform 1 0 25200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_399
timestamp 1663859327
transform 1 0 33152 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_400
timestamp 1663859327
transform 1 0 41104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_401
timestamp 1663859327
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_402
timestamp 1663859327
transform 1 0 13216 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_403
timestamp 1663859327
transform 1 0 21168 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_404
timestamp 1663859327
transform 1 0 29120 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_405
timestamp 1663859327
transform 1 0 37072 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_406
timestamp 1663859327
transform 1 0 45024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_407
timestamp 1663859327
transform 1 0 9296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_408
timestamp 1663859327
transform 1 0 17248 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_409
timestamp 1663859327
transform 1 0 25200 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_410
timestamp 1663859327
transform 1 0 33152 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_411
timestamp 1663859327
transform 1 0 41104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_412
timestamp 1663859327
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_413
timestamp 1663859327
transform 1 0 9184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_414
timestamp 1663859327
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_415
timestamp 1663859327
transform 1 0 17024 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_416
timestamp 1663859327
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_417
timestamp 1663859327
transform 1 0 24864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_418
timestamp 1663859327
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_419
timestamp 1663859327
transform 1 0 32704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_420
timestamp 1663859327
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_421
timestamp 1663859327
transform 1 0 40544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_422
timestamp 1663859327
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _154_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 22512 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _155_
timestamp 1663859327
transform 1 0 13664 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _156_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 21504 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor3_1  _157_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 28112 0 -1 37632
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _158_
timestamp 1663859327
transform -1 0 25984 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _159_
timestamp 1663859327
transform -1 0 36064 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _160_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 17584 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _161_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 32928 0 -1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _162_
timestamp 1663859327
transform 1 0 17584 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _163_
timestamp 1663859327
transform -1 0 26096 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _164_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 22624 0 1 31360
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _165_
timestamp 1663859327
transform -1 0 30800 0 1 42336
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _166_
timestamp 1663859327
transform -1 0 32928 0 -1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _167_
timestamp 1663859327
transform 1 0 11536 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _168_
timestamp 1663859327
transform -1 0 20384 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _169_
timestamp 1663859327
transform -1 0 18704 0 -1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _170_
timestamp 1663859327
transform -1 0 17136 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _171_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 24752 0 -1 40768
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _172_
timestamp 1663859327
transform -1 0 8064 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _173_
timestamp 1663859327
transform -1 0 13104 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _174_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 34384 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _175_
timestamp 1663859327
transform 1 0 12320 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _176_
timestamp 1663859327
transform -1 0 33264 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _177_
timestamp 1663859327
transform 1 0 13104 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _178_
timestamp 1663859327
transform 1 0 8288 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _179_
timestamp 1663859327
transform -1 0 18816 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _180_
timestamp 1663859327
transform -1 0 27888 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _181_
timestamp 1663859327
transform -1 0 10864 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _182_
timestamp 1663859327
transform 1 0 10192 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _183_
timestamp 1663859327
transform 1 0 34272 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1663859327
transform -1 0 36960 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _185_
timestamp 1663859327
transform -1 0 31472 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _186_
timestamp 1663859327
transform -1 0 25088 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _187_
timestamp 1663859327
transform 1 0 29456 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _188_
timestamp 1663859327
transform -1 0 35280 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _189_
timestamp 1663859327
transform -1 0 27216 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _190_
timestamp 1663859327
transform 1 0 8064 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _191_
timestamp 1663859327
transform 1 0 7392 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _192_
timestamp 1663859327
transform 1 0 14560 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _193_
timestamp 1663859327
transform -1 0 13664 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _194_
timestamp 1663859327
transform 1 0 10192 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _195_
timestamp 1663859327
transform -1 0 33264 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _196_
timestamp 1663859327
transform -1 0 11648 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _197_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 11424 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _198_
timestamp 1663859327
transform 1 0 11984 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _199_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 16576 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _200_
timestamp 1663859327
transform -1 0 24192 0 1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _201_
timestamp 1663859327
transform -1 0 22288 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _202_
timestamp 1663859327
transform 1 0 6496 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  _203_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 18704 0 -1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _204_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 12432 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_2  _205_
timestamp 1663859327
transform 1 0 16576 0 1 40768
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__mux4_1  _206_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 21616 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _207_
timestamp 1663859327
transform 1 0 8736 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _208_
timestamp 1663859327
transform -1 0 31248 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _209_
timestamp 1663859327
transform -1 0 22176 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _210_
timestamp 1663859327
transform 1 0 19040 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _211_
timestamp 1663859327
transform -1 0 34384 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _212_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 17584 0 1 34496
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _213_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 11760 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _214_
timestamp 1663859327
transform -1 0 21056 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _215_
timestamp 1663859327
transform -1 0 28672 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _216_
timestamp 1663859327
transform -1 0 32368 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _217_
timestamp 1663859327
transform -1 0 14112 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _218_
timestamp 1663859327
transform -1 0 25088 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _219_
timestamp 1663859327
transform -1 0 34160 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _220_
timestamp 1663859327
transform -1 0 7168 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _221_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 18144 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _222_
timestamp 1663859327
transform 1 0 7840 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _223_
timestamp 1663859327
transform 1 0 11088 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _224_
timestamp 1663859327
transform -1 0 6272 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _225_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 12208 0 -1 39200
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_2  _226_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 31584 0 -1 42336
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _227_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 18480 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _228_
timestamp 1663859327
transform 1 0 13552 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_2  _229_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 24752 0 -1 37632
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _230_
timestamp 1663859327
transform -1 0 8064 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _231_
timestamp 1663859327
transform 1 0 17136 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _232_
timestamp 1663859327
transform 1 0 11872 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _233_
timestamp 1663859327
transform 1 0 13552 0 1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _234_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 27216 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _235_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 19936 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _236_
timestamp 1663859327
transform -1 0 34160 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _237_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 9968 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _238_
timestamp 1663859327
transform -1 0 18928 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _239_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 29456 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _240_
timestamp 1663859327
transform -1 0 29792 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _241_
timestamp 1663859327
transform -1 0 28112 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _242_
timestamp 1663859327
transform -1 0 21056 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _243_
timestamp 1663859327
transform -1 0 31472 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _244_
timestamp 1663859327
transform 1 0 11088 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _245_
timestamp 1663859327
transform 1 0 15456 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _246_
timestamp 1663859327
transform 1 0 28448 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _247_
timestamp 1663859327
transform -1 0 21168 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _248_
timestamp 1663859327
transform -1 0 10192 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _249_
timestamp 1663859327
transform -1 0 7168 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _250_
timestamp 1663859327
transform -1 0 16912 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _251_
timestamp 1663859327
transform 1 0 25536 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _252_
timestamp 1663859327
transform 1 0 28448 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _253_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 32144 0 1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _254_
timestamp 1663859327
transform 1 0 13552 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _255_
timestamp 1663859327
transform 1 0 23408 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _256_
timestamp 1663859327
transform 1 0 28112 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _257_
timestamp 1663859327
transform 1 0 24416 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _258_
timestamp 1663859327
transform 1 0 28336 0 -1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _259_
timestamp 1663859327
transform -1 0 27776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_2  _260_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 24752 0 -1 42336
box -86 -86 2214 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _261_
timestamp 1663859327
transform -1 0 28560 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _262_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 28112 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _263_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 17696 0 -1 37632
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _264_
timestamp 1663859327
transform 1 0 21504 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _265_
timestamp 1663859327
transform -1 0 15792 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _266_
timestamp 1663859327
transform 1 0 14000 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _267_
timestamp 1663859327
transform -1 0 16240 0 1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _268_
timestamp 1663859327
transform 1 0 19376 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _269_
timestamp 1663859327
transform -1 0 35280 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _270_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 31472 0 -1 43904
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _271_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 22960 0 -1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _272_
timestamp 1663859327
transform 1 0 22400 0 -1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _273_
timestamp 1663859327
transform 1 0 31696 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _274_
timestamp 1663859327
transform 1 0 28448 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _275_
timestamp 1663859327
transform 1 0 24080 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _276_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 31584 0 -1 40768
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _277_
timestamp 1663859327
transform -1 0 30576 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _278_
timestamp 1663859327
transform -1 0 30128 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _279_
timestamp 1663859327
transform -1 0 9184 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _280_
timestamp 1663859327
transform 1 0 13552 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _281_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 20608 0 -1 32928
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _282_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 16016 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _283_
timestamp 1663859327
transform -1 0 10192 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _284_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 26656 0 1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _285_
timestamp 1663859327
transform 1 0 11872 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _286_
timestamp 1663859327
transform 1 0 30576 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _287_
timestamp 1663859327
transform 1 0 31696 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _288_
timestamp 1663859327
transform -1 0 29456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _289_
timestamp 1663859327
transform -1 0 19264 0 -1 43904
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _290_
timestamp 1663859327
transform -1 0 32480 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _291_
timestamp 1663859327
transform 1 0 29456 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _292_
timestamp 1663859327
transform -1 0 34832 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _293_
timestamp 1663859327
transform 1 0 14560 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _294_
timestamp 1663859327
transform -1 0 29008 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _295_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 28000 0 1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _296_
timestamp 1663859327
transform -1 0 11984 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _297_
timestamp 1663859327
transform 1 0 29680 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _298_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 16352 0 1 40768
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _299_
timestamp 1663859327
transform 1 0 8960 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _300_
timestamp 1663859327
transform 1 0 25536 0 -1 36064
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _301_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 30240 0 -1 43904
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _302_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 22848 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _303_
timestamp 1663859327
transform -1 0 13664 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _304_
timestamp 1663859327
transform -1 0 24416 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _305_
timestamp 1663859327
transform -1 0 13104 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _306_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 30352 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _307_
timestamp 1663859327
transform 1 0 26208 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _308_
timestamp 1663859327
transform 1 0 28784 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_2  _309_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 26544 0 1 40768
box -86 -86 1990 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _310_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 21504 0 1 40768
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _311_
timestamp 1663859327
transform 1 0 32928 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _312_
timestamp 1663859327
transform 1 0 12208 0 -1 43904
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _313_
timestamp 1663859327
transform -1 0 24304 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _314_
timestamp 1663859327
transform 1 0 10304 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _315_
timestamp 1663859327
transform 1 0 31024 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _316_
timestamp 1663859327
transform 1 0 24976 0 1 36064
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _317_
timestamp 1663859327
transform 1 0 30800 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _318_
timestamp 1663859327
transform -1 0 28784 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _319_
timestamp 1663859327
transform -1 0 9632 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _320_
timestamp 1663859327
transform 1 0 25200 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _321_
timestamp 1663859327
transform -1 0 27104 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _322_
timestamp 1663859327
transform 1 0 22064 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _323_
timestamp 1663859327
transform -1 0 20608 0 1 32928
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _324_
timestamp 1663859327
transform 1 0 10976 0 -1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _325_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 28224 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _326_
timestamp 1663859327
transform 1 0 21840 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _327_
timestamp 1663859327
transform 1 0 19376 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _328_
timestamp 1663859327
transform -1 0 17584 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _329_
timestamp 1663859327
transform 1 0 17808 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _330_
timestamp 1663859327
transform 1 0 13888 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _331_
timestamp 1663859327
transform 1 0 19488 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _332_
timestamp 1663859327
transform 1 0 17808 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _333_
timestamp 1663859327
transform 1 0 13888 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _334_
timestamp 1663859327
transform 1 0 21504 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _335_
timestamp 1663859327
transform 1 0 17808 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _336_
timestamp 1663859327
transform -1 0 22624 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _337_
timestamp 1663859327
transform 1 0 18928 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _338_
timestamp 1663859327
transform 1 0 14336 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _339_
timestamp 1663859327
transform -1 0 28784 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _340_
timestamp 1663859327
transform 1 0 13888 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _341_
timestamp 1663859327
transform -1 0 21056 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _342_
timestamp 1663859327
transform 1 0 17808 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _343_
timestamp 1663859327
transform 1 0 25536 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _344_
timestamp 1663859327
transform 1 0 14336 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _345_
timestamp 1663859327
transform -1 0 21056 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _346_
timestamp 1663859327
transform -1 0 20832 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _347_
timestamp 1663859327
transform -1 0 28784 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _348_
timestamp 1663859327
transform -1 0 24752 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _349_
timestamp 1663859327
transform 1 0 13888 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _350_
timestamp 1663859327
transform 1 0 14336 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _351_
timestamp 1663859327
transform -1 0 13104 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _352_
timestamp 1663859327
transform 1 0 9856 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _353_
timestamp 1663859327
transform -1 0 24752 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _354_
timestamp 1663859327
transform 1 0 14336 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _355_
timestamp 1663859327
transform -1 0 17136 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _356_
timestamp 1663859327
transform -1 0 32704 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _357_
timestamp 1663859327
transform 1 0 10416 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _358_
timestamp 1663859327
transform -1 0 24752 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _359_
timestamp 1663859327
transform 1 0 25536 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _360_
timestamp 1663859327
transform 1 0 24976 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _361_
timestamp 1663859327
transform -1 0 28224 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _362_
timestamp 1663859327
transform 1 0 24976 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _363_
timestamp 1663859327
transform 1 0 10416 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _364_
timestamp 1663859327
transform 1 0 13888 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _365_
timestamp 1663859327
transform -1 0 13104 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _366_ pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 22400 0 -1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _367_
timestamp 1663859327
transform 1 0 19152 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _368_
timestamp 1663859327
transform 1 0 21280 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _369_
timestamp 1663859327
transform 1 0 21504 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _370_
timestamp 1663859327
transform 1 0 21504 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _440_
timestamp 1663859327
transform -1 0 4928 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _441_
timestamp 1663859327
transform -1 0 9296 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  input1 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform 1 0 13440 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1663859327
transform -1 0 48272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1663859327
transform -1 0 48272 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1663859327
transform -1 0 37744 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1663859327
transform 1 0 12208 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1663859327
transform 1 0 1680 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1663859327
transform 1 0 18928 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1663859327
transform -1 0 31696 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output9 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 5152 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output10
timestamp 1663859327
transform 1 0 17584 0 -1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output11
timestamp 1663859327
transform -1 0 36512 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output12
timestamp 1663859327
transform -1 0 3248 0 1 43904
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output13
timestamp 1663859327
transform -1 0 3248 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output14
timestamp 1663859327
transform -1 0 3248 0 1 3136
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output15
timestamp 1663859327
transform -1 0 34608 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_16 pdk/gf180mcuC/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1663859327
transform -1 0 2128 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_17
timestamp 1663859327
transform 1 0 47824 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_18
timestamp 1663859327
transform -1 0 2128 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_19
timestamp 1663859327
transform -1 0 7952 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_20
timestamp 1663859327
transform -1 0 2128 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_21
timestamp 1663859327
transform -1 0 2128 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_22
timestamp 1663859327
transform -1 0 32144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_23
timestamp 1663859327
transform 1 0 47824 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_24
timestamp 1663859327
transform -1 0 38192 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_25
timestamp 1663859327
transform -1 0 3024 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_26
timestamp 1663859327
transform 1 0 8624 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_27
timestamp 1663859327
transform -1 0 35504 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_28
timestamp 1663859327
transform -1 0 2128 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_29
timestamp 1663859327
transform -1 0 2128 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_30
timestamp 1663859327
transform 1 0 47824 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_31
timestamp 1663859327
transform -1 0 2128 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_32
timestamp 1663859327
transform -1 0 2128 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_33
timestamp 1663859327
transform 1 0 47824 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_34
timestamp 1663859327
transform 1 0 47824 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_35
timestamp 1663859327
transform -1 0 42896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_36
timestamp 1663859327
transform 1 0 47824 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_37
timestamp 1663859327
transform -1 0 2800 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_38
timestamp 1663859327
transform -1 0 2128 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_39
timestamp 1663859327
transform -1 0 26768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_40
timestamp 1663859327
transform -1 0 2800 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_41
timestamp 1663859327
transform -1 0 43568 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_42
timestamp 1663859327
transform -1 0 23408 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_43
timestamp 1663859327
transform 1 0 47824 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_44
timestamp 1663859327
transform -1 0 3472 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_45
timestamp 1663859327
transform -1 0 2128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_46
timestamp 1663859327
transform -1 0 9968 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_47
timestamp 1663859327
transform -1 0 18032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_48
timestamp 1663859327
transform -1 0 2128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_49
timestamp 1663859327
transform 1 0 47824 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_50
timestamp 1663859327
transform -1 0 29568 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_51
timestamp 1663859327
transform -1 0 40208 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_52
timestamp 1663859327
transform -1 0 16016 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_53
timestamp 1663859327
transform -1 0 30464 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_54
timestamp 1663859327
transform -1 0 41328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_55
timestamp 1663859327
transform -1 0 2128 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_56
timestamp 1663859327
transform -1 0 6048 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_57
timestamp 1663859327
transform -1 0 2128 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_58
timestamp 1663859327
transform 1 0 46928 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_59
timestamp 1663859327
transform 1 0 47824 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_60
timestamp 1663859327
transform 1 0 47824 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_61
timestamp 1663859327
transform -1 0 38864 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_62
timestamp 1663859327
transform -1 0 2128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_63
timestamp 1663859327
transform 1 0 47824 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_64
timestamp 1663859327
transform -1 0 2128 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_65
timestamp 1663859327
transform -1 0 2128 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_66
timestamp 1663859327
transform 1 0 47824 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_67
timestamp 1663859327
transform -1 0 44240 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_68
timestamp 1663859327
transform -1 0 2128 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_69
timestamp 1663859327
transform 1 0 47824 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_70
timestamp 1663859327
transform -1 0 32368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_71
timestamp 1663859327
transform 1 0 10080 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_72
timestamp 1663859327
transform 1 0 10752 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_73
timestamp 1663859327
transform -1 0 14672 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_74
timestamp 1663859327
transform 1 0 47824 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_75
timestamp 1663859327
transform 1 0 47824 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_76
timestamp 1663859327
transform 1 0 47824 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_77
timestamp 1663859327
transform -1 0 3920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_78
timestamp 1663859327
transform -1 0 46256 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_79
timestamp 1663859327
transform 1 0 47824 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_80
timestamp 1663859327
transform -1 0 2128 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_81
timestamp 1663859327
transform -1 0 2128 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_82
timestamp 1663859327
transform -1 0 21728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_83
timestamp 1663859327
transform 1 0 47824 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  tiny_user_project_84
timestamp 1663859327
transform 1 0 47824 0 1 37632
box -86 -86 534 870
<< labels >>
flabel metal2 s 23520 49200 23632 49800 0 FreeSans 448 90 0 0 io_in[0]
port 0 nsew signal input
flabel metal2 s 49728 49200 49840 49800 0 FreeSans 448 90 0 0 io_in[10]
port 1 nsew signal input
flabel metal2 s 24192 200 24304 800 0 FreeSans 448 90 0 0 io_in[11]
port 2 nsew signal input
flabel metal2 s 11424 49200 11536 49800 0 FreeSans 448 90 0 0 io_in[12]
port 3 nsew signal input
flabel metal2 s 49056 200 49168 800 0 FreeSans 448 90 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 49200 43008 49800 43120 0 FreeSans 448 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 36960 200 37072 800 0 FreeSans 448 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 12096 200 12208 800 0 FreeSans 448 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal3 s 200 47712 800 47824 0 FreeSans 448 0 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 18816 200 18928 800 0 FreeSans 448 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 30912 49200 31024 49800 0 FreeSans 448 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 200 1344 800 1456 0 FreeSans 448 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 33600 200 33712 800 0 FreeSans 448 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal3 s 200 31584 800 31696 0 FreeSans 448 0 0 0 io_in[21]
port 13 nsew signal input
flabel metal3 s 49200 20160 49800 20272 0 FreeSans 448 0 0 0 io_in[22]
port 14 nsew signal input
flabel metal3 s 49200 46368 49800 46480 0 FreeSans 448 0 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s 200 4704 800 4816 0 FreeSans 448 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal2 s 40992 49200 41104 49800 0 FreeSans 448 90 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s 200 40320 800 40432 0 FreeSans 448 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s 49200 14784 49800 14896 0 FreeSans 448 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s 49200 40992 49800 41104 0 FreeSans 448 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal2 s 47712 200 47824 800 0 FreeSans 448 90 0 0 io_in[29]
port 21 nsew signal input
flabel metal2 s 29568 200 29680 800 0 FreeSans 448 90 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s 49200 4032 49800 4144 0 FreeSans 448 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal2 s 14784 49200 14896 49800 0 FreeSans 448 90 0 0 io_in[31]
port 24 nsew signal input
flabel metal2 s 10080 200 10192 800 0 FreeSans 448 90 0 0 io_in[32]
port 25 nsew signal input
flabel metal2 s 25536 49200 25648 49800 0 FreeSans 448 90 0 0 io_in[33]
port 26 nsew signal input
flabel metal2 s 46368 49200 46480 49800 0 FreeSans 448 90 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s 200 12096 800 12208 0 FreeSans 448 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal2 s 16128 49200 16240 49800 0 FreeSans 448 90 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s 49200 45024 49800 45136 0 FreeSans 448 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 49200 25536 49800 25648 0 FreeSans 448 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal2 s 28896 49200 29008 49800 0 FreeSans 448 90 0 0 io_in[4]
port 32 nsew signal input
flabel metal2 s 6720 200 6832 800 0 FreeSans 448 90 0 0 io_in[5]
port 33 nsew signal input
flabel metal2 s 45024 49200 45136 49800 0 FreeSans 448 90 0 0 io_in[6]
port 34 nsew signal input
flabel metal2 s 34272 49200 34384 49800 0 FreeSans 448 90 0 0 io_in[7]
port 35 nsew signal input
flabel metal2 s 6048 49200 6160 49800 0 FreeSans 448 90 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 49200 48384 49800 48496 0 FreeSans 448 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal2 s 15456 200 15568 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 200 8736 800 8848 0 FreeSans 448 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 49200 34272 49800 34384 0 FreeSans 448 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 200 34944 800 35056 0 FreeSans 448 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 200 18816 800 18928 0 FreeSans 448 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 49200 11424 49800 11536 0 FreeSans 448 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 43680 200 43792 800 0 FreeSans 448 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal3 s 200 24192 800 24304 0 FreeSans 448 0 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal3 s 49200 26880 49800 26992 0 FreeSans 448 0 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 21504 49200 21616 49800 0 FreeSans 448 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 12768 49200 12880 49800 0 FreeSans 448 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal2 s 26880 49200 26992 49800 0 FreeSans 448 90 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 18144 49200 18256 49800 0 FreeSans 448 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 14112 200 14224 800 0 FreeSans 448 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal3 s 49200 12768 49800 12880 0 FreeSans 448 0 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal3 s 49200 6048 49800 6160 0 FreeSans 448 0 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s 49200 32256 49800 32368 0 FreeSans 448 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal2 s 3360 200 3472 800 0 FreeSans 448 90 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal2 s 45696 200 45808 800 0 FreeSans 448 90 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s 49200 9408 49800 9520 0 FreeSans 448 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s 200 29568 800 29680 0 FreeSans 448 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s 200 3360 800 3472 0 FreeSans 448 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal2 s 40320 200 40432 800 0 FreeSans 448 90 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal2 s 20832 200 20944 800 0 FreeSans 448 90 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s 49200 16800 49800 16912 0 FreeSans 448 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s 49200 37632 49800 37744 0 FreeSans 448 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s 200 38304 800 38416 0 FreeSans 448 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s 49200 2016 49800 2128 0 FreeSans 448 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s 200 45696 800 45808 0 FreeSans 448 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal2 s 7392 49200 7504 49800 0 FreeSans 448 90 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s 200 32928 800 33040 0 FreeSans 448 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 200 6720 800 6832 0 FreeSans 448 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal2 s 4704 200 4816 800 0 FreeSans 448 90 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 200 20832 800 20944 0 FreeSans 448 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 49200 672 49800 784 0 FreeSans 448 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 49200 28896 49800 29008 0 FreeSans 448 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 49200 18144 49800 18256 0 FreeSans 448 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal2 s 38304 200 38416 800 0 FreeSans 448 90 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 200 36960 800 37072 0 FreeSans 448 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 200 28224 800 28336 0 FreeSans 448 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 200 26208 800 26320 0 FreeSans 448 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 49200 21504 49800 21616 0 FreeSans 448 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 49200 35616 49800 35728 0 FreeSans 448 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal2 s 42336 200 42448 800 0 FreeSans 448 90 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal3 s 49200 39648 49800 39760 0 FreeSans 448 0 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 672 49200 784 49800 0 FreeSans 448 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal3 s 200 10080 800 10192 0 FreeSans 448 0 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 26208 200 26320 800 0 FreeSans 448 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 0 200 112 800 0 FreeSans 448 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal2 s 31584 200 31696 800 0 FreeSans 448 90 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 4032 49200 4144 49800 0 FreeSans 448 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 20160 49200 20272 49800 0 FreeSans 448 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 35616 49200 35728 49800 0 FreeSans 448 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal3 s 200 43680 800 43792 0 FreeSans 448 0 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s 200 22848 800 22960 0 FreeSans 448 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal2 s 1344 200 1456 800 0 FreeSans 448 90 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal2 s 43008 49200 43120 49800 0 FreeSans 448 90 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal2 s 32256 49200 32368 49800 0 FreeSans 448 90 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal2 s 22848 200 22960 800 0 FreeSans 448 90 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal2 s 48384 49200 48496 49800 0 FreeSans 448 90 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 49200 7392 49800 7504 0 FreeSans 448 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s 200 49056 800 49168 0 FreeSans 448 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s 200 17472 800 17584 0 FreeSans 448 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal2 s 8736 200 8848 800 0 FreeSans 448 90 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal2 s 17472 200 17584 800 0 FreeSans 448 90 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s 200 15456 800 15568 0 FreeSans 448 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s 49200 30912 49800 31024 0 FreeSans 448 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal2 s 28224 200 28336 800 0 FreeSans 448 90 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal2 s 39648 49200 39760 49800 0 FreeSans 448 90 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal2 s 37632 49200 37744 49800 0 FreeSans 448 90 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal2 s 2016 49200 2128 49800 0 FreeSans 448 90 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal2 s 9408 49200 9520 49800 0 FreeSans 448 90 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal2 s 34944 200 35056 800 0 FreeSans 448 90 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 200 14112 800 14224 0 FreeSans 448 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 200 42336 800 42448 0 FreeSans 448 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 49200 23520 49800 23632 0 FreeSans 448 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vccd1
port 114 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vssd1
port 115 nsew ground bidirectional
rlabel metal1 24976 46256 24976 46256 0 vccd1
rlabel metal1 24976 45472 24976 45472 0 vssd1
rlabel metal3 35840 41160 35840 41160 0 _000_
rlabel metal2 24920 32704 24920 32704 0 _001_
rlabel metal3 32984 39816 32984 39816 0 _002_
rlabel metal2 26488 30296 26488 30296 0 _003_
rlabel metal2 8232 40936 8232 40936 0 _004_
rlabel metal2 10472 43988 10472 43988 0 _005_
rlabel metal3 11424 45080 11424 45080 0 _006_
rlabel metal3 13440 32760 13440 32760 0 _007_
rlabel metal2 15624 32256 15624 32256 0 _008_
rlabel metal2 17080 33040 17080 33040 0 _009_
rlabel metal2 21952 30968 21952 30968 0 _010_
rlabel metal2 21560 29288 21560 29288 0 _011_
rlabel metal2 19992 39872 19992 39872 0 _012_
rlabel metal3 23352 42392 23352 42392 0 _013_
rlabel metal2 7000 40320 7000 40320 0 _014_
rlabel metal2 4200 39312 4200 39312 0 _015_
rlabel metal4 26264 32648 26264 32648 0 _016_
rlabel metal3 29120 24584 29120 24584 0 _017_
rlabel metal2 4256 44408 4256 44408 0 _018_
rlabel metal3 7952 39368 7952 39368 0 _019_
rlabel metal3 34328 40936 34328 40936 0 _020_
rlabel metal2 15848 35000 15848 35000 0 _021_
rlabel metal2 5152 39368 5152 39368 0 _022_
rlabel metal2 7896 40208 7896 40208 0 _023_
rlabel metal2 3304 46368 3304 46368 0 _024_
rlabel metal2 5880 39088 5880 39088 0 _025_
rlabel metal2 4648 42448 4648 42448 0 _026_
rlabel metal2 24752 35560 24752 35560 0 _027_
rlabel metal2 26152 49112 26152 49112 0 _028_
rlabel metal2 8008 39088 8008 39088 0 _029_
rlabel metal2 19320 39228 19320 39228 0 _030_
rlabel metal4 8008 46648 8008 46648 0 _031_
rlabel metal2 11816 44968 11816 44968 0 _032_
rlabel metal2 5768 39872 5768 39872 0 _033_
rlabel metal3 13328 38696 13328 38696 0 _034_
rlabel metal4 8344 47320 8344 47320 0 _035_
rlabel metal2 5544 43344 5544 43344 0 _036_
rlabel metal3 23128 47376 23128 47376 0 _037_
rlabel metal2 10696 47488 10696 47488 0 _038_
rlabel metal2 21000 32368 21000 32368 0 _039_
rlabel metal2 2744 39592 2744 39592 0 _040_
rlabel metal2 4760 38696 4760 38696 0 _041_
rlabel metal2 26600 47152 26600 47152 0 _042_
rlabel metal2 29568 39816 29568 39816 0 _043_
rlabel metal2 20888 31416 20888 31416 0 _044_
rlabel metal2 30352 39592 30352 39592 0 _045_
rlabel metal3 17416 31640 17416 31640 0 _046_
rlabel metal2 18648 34832 18648 34832 0 _047_
rlabel metal2 30856 41328 30856 41328 0 _048_
rlabel metal2 8120 46984 8120 46984 0 _049_
rlabel metal2 21224 29736 21224 29736 0 _050_
rlabel metal2 20552 29904 20552 29904 0 _051_
rlabel metal2 10920 44072 10920 44072 0 _052_
rlabel metal3 24192 49000 24192 49000 0 _053_
rlabel metal2 15960 34496 15960 34496 0 _054_
rlabel metal2 38920 46928 38920 46928 0 _055_
rlabel metal3 10416 42056 10416 42056 0 _056_
rlabel metal3 7168 41048 7168 41048 0 _057_
rlabel metal3 7448 47096 7448 47096 0 _058_
rlabel metal2 5152 44408 5152 44408 0 _059_
rlabel metal2 26824 31360 26824 31360 0 _060_
rlabel metal4 26768 40040 26768 40040 0 _061_
rlabel metal2 5992 47096 5992 47096 0 _062_
rlabel metal2 21224 44156 21224 44156 0 _063_
rlabel metal3 24808 49336 24808 49336 0 _064_
rlabel metal2 9912 40432 9912 40432 0 _065_
rlabel metal4 24920 33488 24920 33488 0 _066_
rlabel metal3 29568 37352 29568 37352 0 _067_
rlabel metal2 24360 40880 24360 40880 0 _068_
rlabel metal2 24472 41832 24472 41832 0 _069_
rlabel metal2 5880 46200 5880 46200 0 _070_
rlabel metal3 12264 44296 12264 44296 0 _071_
rlabel metal2 21952 39032 21952 39032 0 _072_
rlabel metal3 28448 13272 28448 13272 0 _073_
rlabel metal3 7560 43624 7560 43624 0 _074_
rlabel metal2 2968 40824 2968 40824 0 _075_
rlabel metal3 19600 16408 19600 16408 0 _076_
rlabel metal2 40488 41776 40488 41776 0 _077_
rlabel metal2 35000 42280 35000 42280 0 _078_
rlabel metal3 27776 43512 27776 43512 0 _079_
rlabel metal2 23576 43008 23576 43008 0 _080_
rlabel metal2 22904 34776 22904 34776 0 _081_
rlabel metal2 3976 39592 3976 39592 0 _082_
rlabel metal2 24920 33768 24920 33768 0 _083_
rlabel metal4 24808 31248 24808 31248 0 _084_
rlabel metal2 40712 46816 40712 46816 0 _085_
rlabel metal2 29904 44296 29904 44296 0 _086_
rlabel metal2 5096 40880 5096 40880 0 _087_
rlabel metal3 9240 41832 9240 41832 0 _088_
rlabel metal2 16520 36792 16520 36792 0 _089_
rlabel metal3 19040 35672 19040 35672 0 _090_
rlabel metal3 28784 36456 28784 36456 0 _091_
rlabel metal3 4704 41832 4704 41832 0 _092_
rlabel metal2 29512 44072 29512 44072 0 _093_
rlabel metal3 22792 24248 22792 24248 0 _094_
rlabel metal2 7336 43288 7336 43288 0 _095_
rlabel metal2 29288 36008 29288 36008 0 _096_
rlabel metal3 13832 47320 13832 47320 0 _097_
rlabel metal4 25816 49168 25816 49168 0 _098_
rlabel metal3 30912 44072 30912 44072 0 _099_
rlabel metal2 26600 35504 26600 35504 0 _100_
rlabel metal2 9352 45416 9352 45416 0 _101_
rlabel metal2 27832 46480 27832 46480 0 _102_
rlabel metal2 28728 44968 28728 44968 0 _103_
rlabel metal4 26936 24640 26936 24640 0 _104_
rlabel metal4 26040 49336 26040 49336 0 _105_
rlabel metal2 26376 36120 26376 36120 0 _106_
rlabel metal2 13272 45192 13272 45192 0 _107_
rlabel metal3 17360 24808 17360 24808 0 _108_
rlabel metal2 26488 38080 26488 38080 0 _109_
rlabel metal3 26488 48608 26488 48608 0 _110_
rlabel metal2 24640 44856 24640 44856 0 _111_
rlabel metal2 21840 41160 21840 41160 0 _112_
rlabel metal2 22680 40712 22680 40712 0 _113_
rlabel metal2 12712 45472 12712 45472 0 _114_
rlabel metal2 26320 33432 26320 33432 0 _115_
rlabel metal4 28280 34160 28280 34160 0 _116_
rlabel metal2 27720 42448 27720 42448 0 _117_
rlabel metal2 24248 41216 24248 41216 0 _118_
rlabel metal4 4872 41328 4872 41328 0 _119_
rlabel metal2 2968 26012 2968 26012 0 _120_
rlabel metal3 14784 40488 14784 40488 0 _121_
rlabel metal2 23464 14000 23464 14000 0 _122_
rlabel metal2 26040 36624 26040 36624 0 _123_
rlabel metal2 26152 36848 26152 36848 0 _124_
rlabel metal2 2856 41496 2856 41496 0 _125_
rlabel metal2 25816 47712 25816 47712 0 _126_
rlabel metal2 26376 42336 26376 42336 0 _127_
rlabel metal3 21224 33432 21224 33432 0 _128_
rlabel metal2 19432 33600 19432 33600 0 _129_
rlabel metal3 21168 40376 21168 40376 0 _130_
rlabel metal2 38696 42392 38696 42392 0 _131_
rlabel metal2 22624 33320 22624 33320 0 _132_
rlabel metal2 25648 33320 25648 33320 0 _133_
rlabel metal2 5544 44800 5544 44800 0 _134_
rlabel metal2 22960 41496 22960 41496 0 _135_
rlabel metal2 23576 31416 23576 31416 0 _136_
rlabel metal2 18368 40600 18368 40600 0 _137_
rlabel metal3 24024 31752 24024 31752 0 _138_
rlabel metal2 22848 31864 22848 31864 0 _139_
rlabel metal2 24584 40544 24584 40544 0 _140_
rlabel metal3 22680 26376 22680 26376 0 _141_
rlabel metal2 3976 41552 3976 41552 0 _142_
rlabel metal2 19376 32648 19376 32648 0 _143_
rlabel metal2 17080 33936 17080 33936 0 _144_
rlabel metal2 24472 40432 24472 40432 0 _145_
rlabel metal2 3752 39872 3752 39872 0 _146_
rlabel metal2 7784 40936 7784 40936 0 _147_
rlabel metal2 2632 38192 2632 38192 0 _148_
rlabel metal2 2632 44716 2632 44716 0 _149_
rlabel metal3 23016 24920 23016 24920 0 _150_
rlabel metal3 17472 31752 17472 31752 0 _151_
rlabel metal2 27272 35896 27272 35896 0 _152_
rlabel metal3 18648 11592 18648 11592 0 _153_
rlabel metal2 1960 44352 1960 44352 0 io_in[12]
rlabel metal3 48608 3416 48608 3416 0 io_in[13]
rlabel metal2 48104 43288 48104 43288 0 io_in[14]
rlabel metal3 36736 3416 36736 3416 0 io_in[15]
rlabel metal2 12040 3416 12040 3416 0 io_in[16]
rlabel metal2 1848 46816 1848 46816 0 io_in[17]
rlabel metal2 18760 3416 18760 3416 0 io_in[18]
rlabel metal2 30968 47530 30968 47530 0 io_in[19]
rlabel metal2 4088 47642 4088 47642 0 io_out[20]
rlabel metal2 20216 47250 20216 47250 0 io_out[21]
rlabel metal2 35672 47642 35672 47642 0 io_out[22]
rlabel metal3 1470 43736 1470 43736 0 io_out[23]
rlabel metal3 1414 22904 1414 22904 0 io_out[24]
rlabel metal2 1400 2142 1400 2142 0 io_out[25]
rlabel metal2 33432 46368 33432 46368 0 io_out[27]
rlabel metal2 4144 44968 4144 44968 0 mod.flipflop1.d
rlabel metal2 17024 44968 17024 44968 0 mod.flipflop1.q
rlabel metal2 25928 47096 25928 47096 0 mod.flipflop10.d
rlabel metal2 22008 32928 22008 32928 0 mod.flipflop11.d
rlabel metal2 25256 41216 25256 41216 0 mod.flipflop11.q
rlabel metal2 10752 44184 10752 44184 0 mod.flipflop12.d
rlabel metal2 8288 45304 8288 45304 0 mod.flipflop12.q
rlabel metal3 18928 36456 18928 36456 0 mod.flipflop13.q
rlabel metal2 7560 40992 7560 40992 0 mod.flipflop14.q
rlabel metal2 26544 41832 26544 41832 0 mod.flipflop15.d
rlabel metal3 29008 48440 29008 48440 0 mod.flipflop16.d
rlabel metal2 5992 42560 5992 42560 0 mod.flipflop17.d
rlabel metal2 15176 36120 15176 36120 0 mod.flipflop18.d
rlabel via2 26488 40824 26488 40824 0 mod.flipflop18.q
rlabel metal4 18760 39060 18760 39060 0 mod.flipflop19.q
rlabel metal3 24528 18424 24528 18424 0 mod.flipflop2.d
rlabel metal3 12096 45640 12096 45640 0 mod.flipflop2.q
rlabel metal3 21280 39704 21280 39704 0 mod.flipflop20.q
rlabel metal2 8680 38920 8680 38920 0 mod.flipflop21.d
rlabel metal3 10808 44408 10808 44408 0 mod.flipflop21.q
rlabel metal2 16968 43344 16968 43344 0 mod.flipflop22.q
rlabel metal2 7224 46312 7224 46312 0 mod.flipflop23.q
rlabel metal3 18424 43176 18424 43176 0 mod.flipflop24.q
rlabel metal2 22008 33880 22008 33880 0 mod.flipflop25.q
rlabel metal3 7000 49280 7000 49280 0 mod.flipflop26.q
rlabel metal2 26096 49560 26096 49560 0 mod.flipflop27.d
rlabel metal2 18032 39816 18032 39816 0 mod.flipflop27.q
rlabel metal2 7392 45192 7392 45192 0 mod.flipflop28.q
rlabel metal2 7672 43960 7672 43960 0 mod.flipflop29.d
rlabel metal2 17864 42000 17864 42000 0 mod.flipflop29.q
rlabel metal2 11144 43960 11144 43960 0 mod.flipflop3.q
rlabel metal3 20944 42840 20944 42840 0 mod.flipflop30.q
rlabel metal2 22624 43400 22624 43400 0 mod.flipflop31.q
rlabel metal3 24640 21672 24640 21672 0 mod.flipflop32.d
rlabel metal2 17024 40264 17024 40264 0 mod.flipflop32.q
rlabel metal3 14560 47096 14560 47096 0 mod.flipflop33.d
rlabel metal2 20888 44912 20888 44912 0 mod.flipflop33.q
rlabel metal2 6216 39816 6216 39816 0 mod.flipflop34.d
rlabel metal2 7784 44324 7784 44324 0 mod.flipflop34.q
rlabel metal2 22512 44968 22512 44968 0 mod.flipflop35.q
rlabel metal4 23016 19992 23016 19992 0 mod.flipflop36.q
rlabel metal3 31192 39480 31192 39480 0 mod.flipflop37.d
rlabel metal2 25144 40040 25144 40040 0 mod.flipflop37.q
rlabel metal2 5096 46704 5096 46704 0 mod.flipflop38.q
rlabel metal2 22232 46144 22232 46144 0 mod.flipflop39.q
rlabel metal2 17416 35896 17416 35896 0 mod.flipflop4.q
rlabel metal3 25256 38920 25256 38920 0 mod.flipflop40.q
rlabel metal2 12992 45640 12992 45640 0 mod.flipflop41.d
rlabel metal2 21448 41776 21448 41776 0 mod.flipflop41.q
rlabel metal2 3248 41272 3248 41272 0 mod.flipflop42.q
rlabel metal2 9968 41272 9968 41272 0 mod.flipflop43.q
rlabel metal3 22232 40712 22232 40712 0 mod.flipflop44.q
rlabel metal2 24976 31192 24976 31192 0 mod.flipflop45.q
rlabel metal3 6552 39312 6552 39312 0 mod.flipflop5.q
rlabel metal2 12936 39760 12936 39760 0 mod.flipflop6.q
rlabel metal2 7168 44408 7168 44408 0 mod.flipflop8.d
rlabel metal2 20216 43344 20216 43344 0 mod.flipflop8.q
rlabel metal2 14784 38920 14784 38920 0 mod.flipflop9.d
rlabel metal2 6272 44072 6272 44072 0 net1
rlabel metal2 7336 44744 7336 44744 0 net10
rlabel metal2 20552 39536 20552 39536 0 net11
rlabel metal2 5656 40992 5656 40992 0 net12
rlabel metal2 3304 23128 3304 23128 0 net13
rlabel metal2 3080 3584 3080 3584 0 net14
rlabel metal2 5544 39480 5544 39480 0 net15
rlabel metal3 1302 38360 1302 38360 0 net16
rlabel metal2 48160 4424 48160 4424 0 net17
rlabel metal2 1792 45304 1792 45304 0 net18
rlabel metal2 7560 45752 7560 45752 0 net19
rlabel metal2 47768 18592 47768 18592 0 net2
rlabel metal3 1302 32984 1302 32984 0 net20
rlabel metal3 1302 37016 1302 37016 0 net21
rlabel metal2 31640 2030 31640 2030 0 net22
rlabel metal2 48104 7728 48104 7728 0 net23
rlabel metal2 37800 45752 37800 45752 0 net24
rlabel metal2 2744 46088 2744 46088 0 net25
rlabel metal2 8904 46088 8904 46088 0 net26
rlabel metal2 35000 2030 35000 2030 0 net27
rlabel metal3 1302 14168 1302 14168 0 net28
rlabel metal3 1302 42392 1302 42392 0 net29
rlabel metal2 47768 44688 47768 44688 0 net3
rlabel metal2 48104 23632 48104 23632 0 net30
rlabel metal3 1302 28280 1302 28280 0 net31
rlabel metal3 1302 26264 1302 26264 0 net32
rlabel metal2 48104 21840 48104 21840 0 net33
rlabel metal2 48104 35952 48104 35952 0 net34
rlabel metal2 42392 2030 42392 2030 0 net35
rlabel metal2 48104 40096 48104 40096 0 net36
rlabel metal2 2520 46312 2520 46312 0 net37
rlabel metal3 1302 10136 1302 10136 0 net38
rlabel metal2 26264 2030 26264 2030 0 net39
rlabel metal4 7896 46536 7896 46536 0 net4
rlabel metal2 56 1526 56 1526 0 net40
rlabel metal2 43176 45752 43176 45752 0 net41
rlabel metal2 22904 2030 22904 2030 0 net42
rlabel metal2 48272 45752 48272 45752 0 net43
rlabel metal2 3192 47208 3192 47208 0 net44
rlabel metal3 1302 17528 1302 17528 0 net45
rlabel metal2 8792 1246 8792 1246 0 net46
rlabel metal2 17528 2030 17528 2030 0 net47
rlabel metal3 1302 15512 1302 15512 0 net48
rlabel metal2 48104 31248 48104 31248 0 net49
rlabel metal3 7392 38696 7392 38696 0 net5
rlabel metal2 28280 2030 28280 2030 0 net50
rlabel metal2 39816 45752 39816 45752 0 net51
rlabel metal2 15512 2030 15512 2030 0 net52
rlabel metal3 28560 45752 28560 45752 0 net53
rlabel metal2 40376 1302 40376 1302 0 net54
rlabel metal3 1302 6776 1302 6776 0 net55
rlabel metal2 4760 2030 4760 2030 0 net56
rlabel metal3 1302 20888 1302 20888 0 net57
rlabel metal2 47208 2016 47208 2016 0 net58
rlabel metal2 48104 29232 48104 29232 0 net59
rlabel metal3 4648 44184 4648 44184 0 net6
rlabel metal3 48104 18368 48104 18368 0 net60
rlabel metal2 38360 2030 38360 2030 0 net61
rlabel metal3 1302 8792 1302 8792 0 net62
rlabel metal2 48104 34496 48104 34496 0 net63
rlabel metal3 1302 35000 1302 35000 0 net64
rlabel metal3 1302 18872 1302 18872 0 net65
rlabel metal2 48104 11872 48104 11872 0 net66
rlabel metal2 43736 2030 43736 2030 0 net67
rlabel metal3 1302 24248 1302 24248 0 net68
rlabel metal3 48104 26880 48104 26880 0 net69
rlabel metal2 19432 7392 19432 7392 0 net7
rlabel metal2 21560 49798 21560 49798 0 net70
rlabel metal2 10360 46032 10360 46032 0 net71
rlabel metal3 14616 45752 14616 45752 0 net72
rlabel metal2 14168 2030 14168 2030 0 net73
rlabel metal3 48706 12824 48706 12824 0 net74
rlabel metal2 48104 6272 48104 6272 0 net75
rlabel metal2 48104 32480 48104 32480 0 net76
rlabel metal2 3416 2030 3416 2030 0 net77
rlabel metal2 45752 2030 45752 2030 0 net78
rlabel metal2 48104 9520 48104 9520 0 net79
rlabel metal3 30632 44968 30632 44968 0 net8
rlabel metal3 1302 29624 1302 29624 0 net80
rlabel metal3 1302 3416 1302 3416 0 net81
rlabel metal2 20888 1246 20888 1246 0 net82
rlabel metal2 48104 17136 48104 17136 0 net83
rlabel metal2 48104 37744 48104 37744 0 net84
rlabel metal2 4928 42056 4928 42056 0 net9
<< properties >>
string FIXED_BBOX 0 0 50000 50000
<< end >>
